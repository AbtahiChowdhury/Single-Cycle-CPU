LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE Chowdhury_Package_UnsignedDivider_Dec7 IS
	COMPONENT Chowdhury_UnsignedDivider_Dec7 IS
		PORT(DIVIDEND,DIVISOR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			  QUOTIENT,REMAINDER : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
	END COMPONENT Chowdhury_UnsignedDivider_Dec7;
END PACKAGE Chowdhury_Package_UnsignedDivider_Dec7;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Chowdhury_UnsignedDivider_Dec7 IS
	PORT(DIVIDEND,DIVISOR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		  QUOTIENT,REMAINDER : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END Chowdhury_UnsignedDivider_Dec7;

ARCHITECTURE Chowdhury_Behaviour OF Chowdhury_UnsignedDivider_Dec7 IS
	
	COMPONENT Chowdhury_1BitDiv_Dec7 IS
		PORT(M,SI,BI,OKI : IN STD_LOGIC;
			  BO,OKO,D,SO : OUT STD_LOGIC);
	END COMPONENT;
	
	SIGNAL Q,R : STD_LOGIC_VECTOR(31 DOWNTO 0) := x"00000000";
	
	TYPE SUB_D IS ARRAY (0 TO 1023) OF STD_LOGIC;
	SIGNAL SUB_DS : SUB_D;
	
	TYPE SUB_BO IS ARRAY (0 TO 1023) OF STD_LOGIC;
	SIGNAL SUB_BOS : SUB_BO;
	
	TYPE SUB_OKO IS ARRAY (0 TO 1023) OF STD_LOGIC;
	SIGNAL SUB_OKOS : SUB_OKO;
	
	TYPE SUB_SO IS ARRAY (0 TO 1023) OF STD_LOGIC;
	SIGNAL SUB_SOS : SUB_SO;
	
	TYPE BON IS ARRAY (0 TO 31) OF STD_LOGIC;
	SIGNAL BONS : BON;
	
BEGIN
	
	BONS(0) <= NOT SUB_BOS(31);
	BONS(1) <= NOT SUB_BOS(63);
	BONS(2) <= NOT SUB_BOS(95);
	BONS(3) <= NOT SUB_BOS(127);
	BONS(4) <= NOT SUB_BOS(159);
	BONS(5) <= NOT SUB_BOS(191);
	BONS(6) <= NOT SUB_BOS(223);
	BONS(7) <= NOT SUB_BOS(255);
	BONS(8) <= NOT SUB_BOS(287);
	BONS(9) <= NOT SUB_BOS(319);
	BONS(10) <= NOT SUB_BOS(351);
	BONS(11) <= NOT SUB_BOS(383);
	BONS(12) <= NOT SUB_BOS(415);
	BONS(13) <= NOT SUB_BOS(447);
	BONS(14) <= NOT SUB_BOS(479);
	BONS(15) <= NOT SUB_BOS(511);
	BONS(16) <= NOT SUB_BOS(543);
	BONS(17) <= NOT SUB_BOS(575);
	BONS(18) <= NOT SUB_BOS(607);
	BONS(19) <= NOT SUB_BOS(639);
	BONS(20) <= NOT SUB_BOS(671);
	BONS(21) <= NOT SUB_BOS(703);
	BONS(22) <= NOT SUB_BOS(735);
	BONS(23) <= NOT SUB_BOS(767);
	BONS(24) <= NOT SUB_BOS(799);
	BONS(25) <= NOT SUB_BOS(831);
	BONS(26) <= NOT SUB_BOS(863);
	BONS(27) <= NOT SUB_BOS(895);
	BONS(28) <= NOT SUB_BOS(927);
	BONS(29) <= NOT SUB_BOS(959);
	BONS(30) <= NOT SUB_BOS(991);
	BONS(31) <= NOT SUB_BOS(1023);

	DIV0: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(31), SI=>DIVISOR(0), BI=>'0', OKI=>SUB_OKOS(1), BO=>SUB_BOS(0), OKO=>SUB_OKOS(0), D=>SUB_DS(0), SO=>SUB_SOS(0));
	DIV1: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(1), BI=>SUB_BOS(0), OKI=>SUB_OKOS(2), BO=>SUB_BOS(1), OKO=>SUB_OKOS(1), D=>SUB_DS(1), SO=>SUB_SOS(1));
	DIV2: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(2), BI=>SUB_BOS(1), OKI=>SUB_OKOS(3), BO=>SUB_BOS(2), OKO=>SUB_OKOS(2), D=>SUB_DS(2), SO=>SUB_SOS(2));
	DIV3: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(3), BI=>SUB_BOS(2), OKI=>SUB_OKOS(4), BO=>SUB_BOS(3), OKO=>SUB_OKOS(3), D=>SUB_DS(3), SO=>SUB_SOS(3));
	DIV4: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(4), BI=>SUB_BOS(3), OKI=>SUB_OKOS(5), BO=>SUB_BOS(4), OKO=>SUB_OKOS(4), D=>SUB_DS(4), SO=>SUB_SOS(4));
	DIV5: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(5), BI=>SUB_BOS(4), OKI=>SUB_OKOS(6), BO=>SUB_BOS(5), OKO=>SUB_OKOS(5), D=>SUB_DS(5), SO=>SUB_SOS(5));
	DIV6: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(6), BI=>SUB_BOS(5), OKI=>SUB_OKOS(7), BO=>SUB_BOS(6), OKO=>SUB_OKOS(6), D=>SUB_DS(6), SO=>SUB_SOS(6));
	DIV7: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(7), BI=>SUB_BOS(6), OKI=>SUB_OKOS(8), BO=>SUB_BOS(7), OKO=>SUB_OKOS(7), D=>SUB_DS(7), SO=>SUB_SOS(7));
	DIV8: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(8), BI=>SUB_BOS(7), OKI=>SUB_OKOS(9), BO=>SUB_BOS(8), OKO=>SUB_OKOS(8), D=>SUB_DS(8), SO=>SUB_SOS(8));
	DIV9: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(9), BI=>SUB_BOS(8), OKI=>SUB_OKOS(10), BO=>SUB_BOS(9), OKO=>SUB_OKOS(9), D=>SUB_DS(9), SO=>SUB_SOS(9));
	DIV10: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(10), BI=>SUB_BOS(9), OKI=>SUB_OKOS(11), BO=>SUB_BOS(10), OKO=>SUB_OKOS(10), D=>SUB_DS(10), SO=>SUB_SOS(10));
	DIV11: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(11), BI=>SUB_BOS(10), OKI=>SUB_OKOS(12), BO=>SUB_BOS(11), OKO=>SUB_OKOS(11), D=>SUB_DS(11), SO=>SUB_SOS(11));
	DIV12: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(12), BI=>SUB_BOS(11), OKI=>SUB_OKOS(13), BO=>SUB_BOS(12), OKO=>SUB_OKOS(12), D=>SUB_DS(12), SO=>SUB_SOS(12));
	DIV13: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(13), BI=>SUB_BOS(12), OKI=>SUB_OKOS(14), BO=>SUB_BOS(13), OKO=>SUB_OKOS(13), D=>SUB_DS(13), SO=>SUB_SOS(13));
	DIV14: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(14), BI=>SUB_BOS(13), OKI=>SUB_OKOS(15), BO=>SUB_BOS(14), OKO=>SUB_OKOS(14), D=>SUB_DS(14), SO=>SUB_SOS(14));
	DIV15: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(15), BI=>SUB_BOS(14), OKI=>SUB_OKOS(16), BO=>SUB_BOS(15), OKO=>SUB_OKOS(15), D=>SUB_DS(15), SO=>SUB_SOS(15));
	DIV16: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(16), BI=>SUB_BOS(15), OKI=>SUB_OKOS(17), BO=>SUB_BOS(16), OKO=>SUB_OKOS(16), D=>SUB_DS(16), SO=>SUB_SOS(16));
	DIV17: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(17), BI=>SUB_BOS(16), OKI=>SUB_OKOS(18), BO=>SUB_BOS(17), OKO=>SUB_OKOS(17), D=>SUB_DS(17), SO=>SUB_SOS(17));
	DIV18: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(18), BI=>SUB_BOS(17), OKI=>SUB_OKOS(19), BO=>SUB_BOS(18), OKO=>SUB_OKOS(18), D=>SUB_DS(18), SO=>SUB_SOS(18));
	DIV19: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(19), BI=>SUB_BOS(18), OKI=>SUB_OKOS(20), BO=>SUB_BOS(19), OKO=>SUB_OKOS(19), D=>SUB_DS(19), SO=>SUB_SOS(19));
	DIV20: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(20), BI=>SUB_BOS(19), OKI=>SUB_OKOS(21), BO=>SUB_BOS(20), OKO=>SUB_OKOS(20), D=>SUB_DS(20), SO=>SUB_SOS(20));
	DIV21: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(21), BI=>SUB_BOS(20), OKI=>SUB_OKOS(22), BO=>SUB_BOS(21), OKO=>SUB_OKOS(21), D=>SUB_DS(21), SO=>SUB_SOS(21));
	DIV22: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(22), BI=>SUB_BOS(21), OKI=>SUB_OKOS(23), BO=>SUB_BOS(22), OKO=>SUB_OKOS(22), D=>SUB_DS(22), SO=>SUB_SOS(22));
	DIV23: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(23), BI=>SUB_BOS(22), OKI=>SUB_OKOS(24), BO=>SUB_BOS(23), OKO=>SUB_OKOS(23), D=>SUB_DS(23), SO=>SUB_SOS(23));
	DIV24: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(24), BI=>SUB_BOS(23), OKI=>SUB_OKOS(25), BO=>SUB_BOS(24), OKO=>SUB_OKOS(24), D=>SUB_DS(24), SO=>SUB_SOS(24));
	DIV25: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(25), BI=>SUB_BOS(24), OKI=>SUB_OKOS(26), BO=>SUB_BOS(25), OKO=>SUB_OKOS(25), D=>SUB_DS(25), SO=>SUB_SOS(25));
	DIV26: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(26), BI=>SUB_BOS(25), OKI=>SUB_OKOS(27), BO=>SUB_BOS(26), OKO=>SUB_OKOS(26), D=>SUB_DS(26), SO=>SUB_SOS(26));
	DIV27: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(27), BI=>SUB_BOS(26), OKI=>SUB_OKOS(28), BO=>SUB_BOS(27), OKO=>SUB_OKOS(27), D=>SUB_DS(27), SO=>SUB_SOS(27));
	DIV28: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(28), BI=>SUB_BOS(27), OKI=>SUB_OKOS(29), BO=>SUB_BOS(28), OKO=>SUB_OKOS(28), D=>SUB_DS(28), SO=>SUB_SOS(28));
	DIV29: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(29), BI=>SUB_BOS(28), OKI=>SUB_OKOS(30), BO=>SUB_BOS(29), OKO=>SUB_OKOS(29), D=>SUB_DS(29), SO=>SUB_SOS(29));
	DIV30: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(30), BI=>SUB_BOS(29), OKI=>SUB_OKOS(31), BO=>SUB_BOS(30), OKO=>SUB_OKOS(30), D=>SUB_DS(30), SO=>SUB_SOS(30));
	DIV31: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>'0', SI=>DIVISOR(31), BI=>SUB_BOS(30), OKI=>BONS(0), BO=>SUB_BOS(31), OKO=>SUB_OKOS(31), D=>SUB_DS(31), SO=>SUB_SOS(31));

	DIV32: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(30), SI=>SUB_SOS(0), BI=>'0', OKI=>SUB_OKOS(33), BO=>SUB_BOS(32), OKO=>SUB_OKOS(32), D=>SUB_DS(32), SO=>SUB_SOS(32));
	DIV33: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(0), SI=>SUB_SOS(1), BI=>SUB_BOS(32), OKI=>SUB_OKOS(34), BO=>SUB_BOS(33), OKO=>SUB_OKOS(33), D=>SUB_DS(33), SO=>SUB_SOS(33));
	DIV34: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(1), SI=>SUB_SOS(2), BI=>SUB_BOS(33), OKI=>SUB_OKOS(35), BO=>SUB_BOS(34), OKO=>SUB_OKOS(34), D=>SUB_DS(34), SO=>SUB_SOS(34));
	DIV35: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(2), SI=>SUB_SOS(3), BI=>SUB_BOS(34), OKI=>SUB_OKOS(36), BO=>SUB_BOS(35), OKO=>SUB_OKOS(35), D=>SUB_DS(35), SO=>SUB_SOS(35));
	DIV36: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(3), SI=>SUB_SOS(4), BI=>SUB_BOS(35), OKI=>SUB_OKOS(37), BO=>SUB_BOS(36), OKO=>SUB_OKOS(36), D=>SUB_DS(36), SO=>SUB_SOS(36));
	DIV37: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(4), SI=>SUB_SOS(5), BI=>SUB_BOS(36), OKI=>SUB_OKOS(38), BO=>SUB_BOS(37), OKO=>SUB_OKOS(37), D=>SUB_DS(37), SO=>SUB_SOS(37));
	DIV38: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(5), SI=>SUB_SOS(6), BI=>SUB_BOS(37), OKI=>SUB_OKOS(39), BO=>SUB_BOS(38), OKO=>SUB_OKOS(38), D=>SUB_DS(38), SO=>SUB_SOS(38));
	DIV39: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(6), SI=>SUB_SOS(7), BI=>SUB_BOS(38), OKI=>SUB_OKOS(40), BO=>SUB_BOS(39), OKO=>SUB_OKOS(39), D=>SUB_DS(39), SO=>SUB_SOS(39));
	DIV40: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(7), SI=>SUB_SOS(8), BI=>SUB_BOS(39), OKI=>SUB_OKOS(41), BO=>SUB_BOS(40), OKO=>SUB_OKOS(40), D=>SUB_DS(40), SO=>SUB_SOS(40));
	DIV41: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(8), SI=>SUB_SOS(9), BI=>SUB_BOS(40), OKI=>SUB_OKOS(42), BO=>SUB_BOS(41), OKO=>SUB_OKOS(41), D=>SUB_DS(41), SO=>SUB_SOS(41));
	DIV42: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(9), SI=>SUB_SOS(10), BI=>SUB_BOS(41), OKI=>SUB_OKOS(43), BO=>SUB_BOS(42), OKO=>SUB_OKOS(42), D=>SUB_DS(42), SO=>SUB_SOS(42));
	DIV43: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(10), SI=>SUB_SOS(11), BI=>SUB_BOS(42), OKI=>SUB_OKOS(44), BO=>SUB_BOS(43), OKO=>SUB_OKOS(43), D=>SUB_DS(43), SO=>SUB_SOS(43));
	DIV44: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(11), SI=>SUB_SOS(12), BI=>SUB_BOS(43), OKI=>SUB_OKOS(45), BO=>SUB_BOS(44), OKO=>SUB_OKOS(44), D=>SUB_DS(44), SO=>SUB_SOS(44));
	DIV45: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(12), SI=>SUB_SOS(13), BI=>SUB_BOS(44), OKI=>SUB_OKOS(46), BO=>SUB_BOS(45), OKO=>SUB_OKOS(45), D=>SUB_DS(45), SO=>SUB_SOS(45));
	DIV46: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(13), SI=>SUB_SOS(14), BI=>SUB_BOS(45), OKI=>SUB_OKOS(47), BO=>SUB_BOS(46), OKO=>SUB_OKOS(46), D=>SUB_DS(46), SO=>SUB_SOS(46));
	DIV47: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(14), SI=>SUB_SOS(15), BI=>SUB_BOS(46), OKI=>SUB_OKOS(48), BO=>SUB_BOS(47), OKO=>SUB_OKOS(47), D=>SUB_DS(47), SO=>SUB_SOS(47));
	DIV48: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(15), SI=>SUB_SOS(16), BI=>SUB_BOS(47), OKI=>SUB_OKOS(49), BO=>SUB_BOS(48), OKO=>SUB_OKOS(48), D=>SUB_DS(48), SO=>SUB_SOS(48));
	DIV49: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(16), SI=>SUB_SOS(17), BI=>SUB_BOS(48), OKI=>SUB_OKOS(50), BO=>SUB_BOS(49), OKO=>SUB_OKOS(49), D=>SUB_DS(49), SO=>SUB_SOS(49));
	DIV50: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(17), SI=>SUB_SOS(18), BI=>SUB_BOS(49), OKI=>SUB_OKOS(51), BO=>SUB_BOS(50), OKO=>SUB_OKOS(50), D=>SUB_DS(50), SO=>SUB_SOS(50));
	DIV51: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(18), SI=>SUB_SOS(19), BI=>SUB_BOS(50), OKI=>SUB_OKOS(52), BO=>SUB_BOS(51), OKO=>SUB_OKOS(51), D=>SUB_DS(51), SO=>SUB_SOS(51));
	DIV52: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(19), SI=>SUB_SOS(20), BI=>SUB_BOS(51), OKI=>SUB_OKOS(53), BO=>SUB_BOS(52), OKO=>SUB_OKOS(52), D=>SUB_DS(52), SO=>SUB_SOS(52));
	DIV53: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(20), SI=>SUB_SOS(21), BI=>SUB_BOS(52), OKI=>SUB_OKOS(54), BO=>SUB_BOS(53), OKO=>SUB_OKOS(53), D=>SUB_DS(53), SO=>SUB_SOS(53));
	DIV54: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(21), SI=>SUB_SOS(22), BI=>SUB_BOS(53), OKI=>SUB_OKOS(55), BO=>SUB_BOS(54), OKO=>SUB_OKOS(54), D=>SUB_DS(54), SO=>SUB_SOS(54));
	DIV55: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(22), SI=>SUB_SOS(23), BI=>SUB_BOS(54), OKI=>SUB_OKOS(56), BO=>SUB_BOS(55), OKO=>SUB_OKOS(55), D=>SUB_DS(55), SO=>SUB_SOS(55));
	DIV56: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(23), SI=>SUB_SOS(24), BI=>SUB_BOS(55), OKI=>SUB_OKOS(57), BO=>SUB_BOS(56), OKO=>SUB_OKOS(56), D=>SUB_DS(56), SO=>SUB_SOS(56));
	DIV57: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(24), SI=>SUB_SOS(25), BI=>SUB_BOS(56), OKI=>SUB_OKOS(58), BO=>SUB_BOS(57), OKO=>SUB_OKOS(57), D=>SUB_DS(57), SO=>SUB_SOS(57));
	DIV58: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(25), SI=>SUB_SOS(26), BI=>SUB_BOS(57), OKI=>SUB_OKOS(59), BO=>SUB_BOS(58), OKO=>SUB_OKOS(58), D=>SUB_DS(58), SO=>SUB_SOS(58));
	DIV59: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(26), SI=>SUB_SOS(27), BI=>SUB_BOS(58), OKI=>SUB_OKOS(60), BO=>SUB_BOS(59), OKO=>SUB_OKOS(59), D=>SUB_DS(59), SO=>SUB_SOS(59));
	DIV60: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(27), SI=>SUB_SOS(28), BI=>SUB_BOS(59), OKI=>SUB_OKOS(61), BO=>SUB_BOS(60), OKO=>SUB_OKOS(60), D=>SUB_DS(60), SO=>SUB_SOS(60));
	DIV61: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(28), SI=>SUB_SOS(29), BI=>SUB_BOS(60), OKI=>SUB_OKOS(62), BO=>SUB_BOS(61), OKO=>SUB_OKOS(61), D=>SUB_DS(61), SO=>SUB_SOS(61));
	DIV62: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(29), SI=>SUB_SOS(30), BI=>SUB_BOS(61), OKI=>SUB_OKOS(63), BO=>SUB_BOS(62), OKO=>SUB_OKOS(62), D=>SUB_DS(62), SO=>SUB_SOS(62));
	DIV63: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(30), SI=>SUB_SOS(31), BI=>SUB_BOS(62), OKI=>BONS(1), BO=>SUB_BOS(63), OKO=>SUB_OKOS(63), D=>SUB_DS(63), SO=>SUB_SOS(63));

	DIV64: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(29), SI=>SUB_SOS(32), BI=>'0', OKI=>SUB_OKOS(65), BO=>SUB_BOS(64), OKO=>SUB_OKOS(64), D=>SUB_DS(64), SO=>SUB_SOS(64));
	DIV65: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(32), SI=>SUB_SOS(33), BI=>SUB_BOS(64), OKI=>SUB_OKOS(66), BO=>SUB_BOS(65), OKO=>SUB_OKOS(65), D=>SUB_DS(65), SO=>SUB_SOS(65));
	DIV66: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(33), SI=>SUB_SOS(34), BI=>SUB_BOS(65), OKI=>SUB_OKOS(67), BO=>SUB_BOS(66), OKO=>SUB_OKOS(66), D=>SUB_DS(66), SO=>SUB_SOS(66));
	DIV67: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(34), SI=>SUB_SOS(35), BI=>SUB_BOS(66), OKI=>SUB_OKOS(68), BO=>SUB_BOS(67), OKO=>SUB_OKOS(67), D=>SUB_DS(67), SO=>SUB_SOS(67));
	DIV68: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(35), SI=>SUB_SOS(36), BI=>SUB_BOS(67), OKI=>SUB_OKOS(69), BO=>SUB_BOS(68), OKO=>SUB_OKOS(68), D=>SUB_DS(68), SO=>SUB_SOS(68));
	DIV69: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(36), SI=>SUB_SOS(37), BI=>SUB_BOS(68), OKI=>SUB_OKOS(70), BO=>SUB_BOS(69), OKO=>SUB_OKOS(69), D=>SUB_DS(69), SO=>SUB_SOS(69));
	DIV70: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(37), SI=>SUB_SOS(38), BI=>SUB_BOS(69), OKI=>SUB_OKOS(71), BO=>SUB_BOS(70), OKO=>SUB_OKOS(70), D=>SUB_DS(70), SO=>SUB_SOS(70));
	DIV71: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(38), SI=>SUB_SOS(39), BI=>SUB_BOS(70), OKI=>SUB_OKOS(72), BO=>SUB_BOS(71), OKO=>SUB_OKOS(71), D=>SUB_DS(71), SO=>SUB_SOS(71));
	DIV72: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(39), SI=>SUB_SOS(40), BI=>SUB_BOS(71), OKI=>SUB_OKOS(73), BO=>SUB_BOS(72), OKO=>SUB_OKOS(72), D=>SUB_DS(72), SO=>SUB_SOS(72));
	DIV73: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(40), SI=>SUB_SOS(41), BI=>SUB_BOS(72), OKI=>SUB_OKOS(74), BO=>SUB_BOS(73), OKO=>SUB_OKOS(73), D=>SUB_DS(73), SO=>SUB_SOS(73));
	DIV74: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(41), SI=>SUB_SOS(42), BI=>SUB_BOS(73), OKI=>SUB_OKOS(75), BO=>SUB_BOS(74), OKO=>SUB_OKOS(74), D=>SUB_DS(74), SO=>SUB_SOS(74));
	DIV75: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(42), SI=>SUB_SOS(43), BI=>SUB_BOS(74), OKI=>SUB_OKOS(76), BO=>SUB_BOS(75), OKO=>SUB_OKOS(75), D=>SUB_DS(75), SO=>SUB_SOS(75));
	DIV76: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(43), SI=>SUB_SOS(44), BI=>SUB_BOS(75), OKI=>SUB_OKOS(77), BO=>SUB_BOS(76), OKO=>SUB_OKOS(76), D=>SUB_DS(76), SO=>SUB_SOS(76));
	DIV77: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(44), SI=>SUB_SOS(45), BI=>SUB_BOS(76), OKI=>SUB_OKOS(78), BO=>SUB_BOS(77), OKO=>SUB_OKOS(77), D=>SUB_DS(77), SO=>SUB_SOS(77));
	DIV78: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(45), SI=>SUB_SOS(46), BI=>SUB_BOS(77), OKI=>SUB_OKOS(79), BO=>SUB_BOS(78), OKO=>SUB_OKOS(78), D=>SUB_DS(78), SO=>SUB_SOS(78));
	DIV79: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(46), SI=>SUB_SOS(47), BI=>SUB_BOS(78), OKI=>SUB_OKOS(80), BO=>SUB_BOS(79), OKO=>SUB_OKOS(79), D=>SUB_DS(79), SO=>SUB_SOS(79));
	DIV80: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(47), SI=>SUB_SOS(48), BI=>SUB_BOS(79), OKI=>SUB_OKOS(81), BO=>SUB_BOS(80), OKO=>SUB_OKOS(80), D=>SUB_DS(80), SO=>SUB_SOS(80));
	DIV81: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(48), SI=>SUB_SOS(49), BI=>SUB_BOS(80), OKI=>SUB_OKOS(82), BO=>SUB_BOS(81), OKO=>SUB_OKOS(81), D=>SUB_DS(81), SO=>SUB_SOS(81));
	DIV82: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(49), SI=>SUB_SOS(50), BI=>SUB_BOS(81), OKI=>SUB_OKOS(83), BO=>SUB_BOS(82), OKO=>SUB_OKOS(82), D=>SUB_DS(82), SO=>SUB_SOS(82));
	DIV83: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(50), SI=>SUB_SOS(51), BI=>SUB_BOS(82), OKI=>SUB_OKOS(84), BO=>SUB_BOS(83), OKO=>SUB_OKOS(83), D=>SUB_DS(83), SO=>SUB_SOS(83));
	DIV84: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(51), SI=>SUB_SOS(52), BI=>SUB_BOS(83), OKI=>SUB_OKOS(85), BO=>SUB_BOS(84), OKO=>SUB_OKOS(84), D=>SUB_DS(84), SO=>SUB_SOS(84));
	DIV85: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(52), SI=>SUB_SOS(53), BI=>SUB_BOS(84), OKI=>SUB_OKOS(86), BO=>SUB_BOS(85), OKO=>SUB_OKOS(85), D=>SUB_DS(85), SO=>SUB_SOS(85));
	DIV86: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(53), SI=>SUB_SOS(54), BI=>SUB_BOS(85), OKI=>SUB_OKOS(87), BO=>SUB_BOS(86), OKO=>SUB_OKOS(86), D=>SUB_DS(86), SO=>SUB_SOS(86));
	DIV87: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(54), SI=>SUB_SOS(55), BI=>SUB_BOS(86), OKI=>SUB_OKOS(88), BO=>SUB_BOS(87), OKO=>SUB_OKOS(87), D=>SUB_DS(87), SO=>SUB_SOS(87));
	DIV88: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(55), SI=>SUB_SOS(56), BI=>SUB_BOS(87), OKI=>SUB_OKOS(89), BO=>SUB_BOS(88), OKO=>SUB_OKOS(88), D=>SUB_DS(88), SO=>SUB_SOS(88));
	DIV89: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(56), SI=>SUB_SOS(57), BI=>SUB_BOS(88), OKI=>SUB_OKOS(90), BO=>SUB_BOS(89), OKO=>SUB_OKOS(89), D=>SUB_DS(89), SO=>SUB_SOS(89));
	DIV90: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(57), SI=>SUB_SOS(58), BI=>SUB_BOS(89), OKI=>SUB_OKOS(91), BO=>SUB_BOS(90), OKO=>SUB_OKOS(90), D=>SUB_DS(90), SO=>SUB_SOS(90));
	DIV91: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(58), SI=>SUB_SOS(59), BI=>SUB_BOS(90), OKI=>SUB_OKOS(92), BO=>SUB_BOS(91), OKO=>SUB_OKOS(91), D=>SUB_DS(91), SO=>SUB_SOS(91));
	DIV92: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(59), SI=>SUB_SOS(60), BI=>SUB_BOS(91), OKI=>SUB_OKOS(93), BO=>SUB_BOS(92), OKO=>SUB_OKOS(92), D=>SUB_DS(92), SO=>SUB_SOS(92));
	DIV93: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(60), SI=>SUB_SOS(61), BI=>SUB_BOS(92), OKI=>SUB_OKOS(94), BO=>SUB_BOS(93), OKO=>SUB_OKOS(93), D=>SUB_DS(93), SO=>SUB_SOS(93));
	DIV94: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(61), SI=>SUB_SOS(62), BI=>SUB_BOS(93), OKI=>SUB_OKOS(95), BO=>SUB_BOS(94), OKO=>SUB_OKOS(94), D=>SUB_DS(94), SO=>SUB_SOS(94));
	DIV95: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(62), SI=>SUB_SOS(63), BI=>SUB_BOS(94), OKI=>BONS(2), BO=>SUB_BOS(95), OKO=>SUB_OKOS(95), D=>SUB_DS(95), SO=>SUB_SOS(95));

	DIV96: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(28), SI=>SUB_SOS(64), BI=>'0', OKI=>SUB_OKOS(97), BO=>SUB_BOS(96), OKO=>SUB_OKOS(96), D=>SUB_DS(96), SO=>SUB_SOS(96));
	DIV97: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(64), SI=>SUB_SOS(65), BI=>SUB_BOS(96), OKI=>SUB_OKOS(98), BO=>SUB_BOS(97), OKO=>SUB_OKOS(97), D=>SUB_DS(97), SO=>SUB_SOS(97));
	DIV98: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(65), SI=>SUB_SOS(66), BI=>SUB_BOS(97), OKI=>SUB_OKOS(99), BO=>SUB_BOS(98), OKO=>SUB_OKOS(98), D=>SUB_DS(98), SO=>SUB_SOS(98));
	DIV99: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(66), SI=>SUB_SOS(67), BI=>SUB_BOS(98), OKI=>SUB_OKOS(100), BO=>SUB_BOS(99), OKO=>SUB_OKOS(99), D=>SUB_DS(99), SO=>SUB_SOS(99));
	DIV100: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(67), SI=>SUB_SOS(68), BI=>SUB_BOS(99), OKI=>SUB_OKOS(101), BO=>SUB_BOS(100), OKO=>SUB_OKOS(100), D=>SUB_DS(100), SO=>SUB_SOS(100));
	DIV101: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(68), SI=>SUB_SOS(69), BI=>SUB_BOS(100), OKI=>SUB_OKOS(102), BO=>SUB_BOS(101), OKO=>SUB_OKOS(101), D=>SUB_DS(101), SO=>SUB_SOS(101));
	DIV102: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(69), SI=>SUB_SOS(70), BI=>SUB_BOS(101), OKI=>SUB_OKOS(103), BO=>SUB_BOS(102), OKO=>SUB_OKOS(102), D=>SUB_DS(102), SO=>SUB_SOS(102));
	DIV103: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(70), SI=>SUB_SOS(71), BI=>SUB_BOS(102), OKI=>SUB_OKOS(104), BO=>SUB_BOS(103), OKO=>SUB_OKOS(103), D=>SUB_DS(103), SO=>SUB_SOS(103));
	DIV104: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(71), SI=>SUB_SOS(72), BI=>SUB_BOS(103), OKI=>SUB_OKOS(105), BO=>SUB_BOS(104), OKO=>SUB_OKOS(104), D=>SUB_DS(104), SO=>SUB_SOS(104));
	DIV105: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(72), SI=>SUB_SOS(73), BI=>SUB_BOS(104), OKI=>SUB_OKOS(106), BO=>SUB_BOS(105), OKO=>SUB_OKOS(105), D=>SUB_DS(105), SO=>SUB_SOS(105));
	DIV106: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(73), SI=>SUB_SOS(74), BI=>SUB_BOS(105), OKI=>SUB_OKOS(107), BO=>SUB_BOS(106), OKO=>SUB_OKOS(106), D=>SUB_DS(106), SO=>SUB_SOS(106));
	DIV107: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(74), SI=>SUB_SOS(75), BI=>SUB_BOS(106), OKI=>SUB_OKOS(108), BO=>SUB_BOS(107), OKO=>SUB_OKOS(107), D=>SUB_DS(107), SO=>SUB_SOS(107));
	DIV108: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(75), SI=>SUB_SOS(76), BI=>SUB_BOS(107), OKI=>SUB_OKOS(109), BO=>SUB_BOS(108), OKO=>SUB_OKOS(108), D=>SUB_DS(108), SO=>SUB_SOS(108));
	DIV109: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(76), SI=>SUB_SOS(77), BI=>SUB_BOS(108), OKI=>SUB_OKOS(110), BO=>SUB_BOS(109), OKO=>SUB_OKOS(109), D=>SUB_DS(109), SO=>SUB_SOS(109));
	DIV110: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(77), SI=>SUB_SOS(78), BI=>SUB_BOS(109), OKI=>SUB_OKOS(111), BO=>SUB_BOS(110), OKO=>SUB_OKOS(110), D=>SUB_DS(110), SO=>SUB_SOS(110));
	DIV111: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(78), SI=>SUB_SOS(79), BI=>SUB_BOS(110), OKI=>SUB_OKOS(112), BO=>SUB_BOS(111), OKO=>SUB_OKOS(111), D=>SUB_DS(111), SO=>SUB_SOS(111));
	DIV112: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(79), SI=>SUB_SOS(80), BI=>SUB_BOS(111), OKI=>SUB_OKOS(113), BO=>SUB_BOS(112), OKO=>SUB_OKOS(112), D=>SUB_DS(112), SO=>SUB_SOS(112));
	DIV113: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(80), SI=>SUB_SOS(81), BI=>SUB_BOS(112), OKI=>SUB_OKOS(114), BO=>SUB_BOS(113), OKO=>SUB_OKOS(113), D=>SUB_DS(113), SO=>SUB_SOS(113));
	DIV114: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(81), SI=>SUB_SOS(82), BI=>SUB_BOS(113), OKI=>SUB_OKOS(115), BO=>SUB_BOS(114), OKO=>SUB_OKOS(114), D=>SUB_DS(114), SO=>SUB_SOS(114));
	DIV115: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(82), SI=>SUB_SOS(83), BI=>SUB_BOS(114), OKI=>SUB_OKOS(116), BO=>SUB_BOS(115), OKO=>SUB_OKOS(115), D=>SUB_DS(115), SO=>SUB_SOS(115));
	DIV116: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(83), SI=>SUB_SOS(84), BI=>SUB_BOS(115), OKI=>SUB_OKOS(117), BO=>SUB_BOS(116), OKO=>SUB_OKOS(116), D=>SUB_DS(116), SO=>SUB_SOS(116));
	DIV117: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(84), SI=>SUB_SOS(85), BI=>SUB_BOS(116), OKI=>SUB_OKOS(118), BO=>SUB_BOS(117), OKO=>SUB_OKOS(117), D=>SUB_DS(117), SO=>SUB_SOS(117));
	DIV118: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(85), SI=>SUB_SOS(86), BI=>SUB_BOS(117), OKI=>SUB_OKOS(119), BO=>SUB_BOS(118), OKO=>SUB_OKOS(118), D=>SUB_DS(118), SO=>SUB_SOS(118));
	DIV119: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(86), SI=>SUB_SOS(87), BI=>SUB_BOS(118), OKI=>SUB_OKOS(120), BO=>SUB_BOS(119), OKO=>SUB_OKOS(119), D=>SUB_DS(119), SO=>SUB_SOS(119));
	DIV120: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(87), SI=>SUB_SOS(88), BI=>SUB_BOS(119), OKI=>SUB_OKOS(121), BO=>SUB_BOS(120), OKO=>SUB_OKOS(120), D=>SUB_DS(120), SO=>SUB_SOS(120));
	DIV121: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(88), SI=>SUB_SOS(89), BI=>SUB_BOS(120), OKI=>SUB_OKOS(122), BO=>SUB_BOS(121), OKO=>SUB_OKOS(121), D=>SUB_DS(121), SO=>SUB_SOS(121));
	DIV122: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(89), SI=>SUB_SOS(90), BI=>SUB_BOS(121), OKI=>SUB_OKOS(123), BO=>SUB_BOS(122), OKO=>SUB_OKOS(122), D=>SUB_DS(122), SO=>SUB_SOS(122));
	DIV123: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(90), SI=>SUB_SOS(91), BI=>SUB_BOS(122), OKI=>SUB_OKOS(124), BO=>SUB_BOS(123), OKO=>SUB_OKOS(123), D=>SUB_DS(123), SO=>SUB_SOS(123));
	DIV124: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(91), SI=>SUB_SOS(92), BI=>SUB_BOS(123), OKI=>SUB_OKOS(125), BO=>SUB_BOS(124), OKO=>SUB_OKOS(124), D=>SUB_DS(124), SO=>SUB_SOS(124));
	DIV125: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(92), SI=>SUB_SOS(93), BI=>SUB_BOS(124), OKI=>SUB_OKOS(126), BO=>SUB_BOS(125), OKO=>SUB_OKOS(125), D=>SUB_DS(125), SO=>SUB_SOS(125));
	DIV126: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(93), SI=>SUB_SOS(94), BI=>SUB_BOS(125), OKI=>SUB_OKOS(127), BO=>SUB_BOS(126), OKO=>SUB_OKOS(126), D=>SUB_DS(126), SO=>SUB_SOS(126));
	DIV127: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(94), SI=>SUB_SOS(95), BI=>SUB_BOS(126), OKI=>BONS(3), BO=>SUB_BOS(127), OKO=>SUB_OKOS(127), D=>SUB_DS(127), SO=>SUB_SOS(127));

	DIV128: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(27), SI=>SUB_SOS(96), BI=>'0', OKI=>SUB_OKOS(129), BO=>SUB_BOS(128), OKO=>SUB_OKOS(128), D=>SUB_DS(128), SO=>SUB_SOS(128));
	DIV129: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(96), SI=>SUB_SOS(97), BI=>SUB_BOS(128), OKI=>SUB_OKOS(130), BO=>SUB_BOS(129), OKO=>SUB_OKOS(129), D=>SUB_DS(129), SO=>SUB_SOS(129));
	DIV130: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(97), SI=>SUB_SOS(98), BI=>SUB_BOS(129), OKI=>SUB_OKOS(131), BO=>SUB_BOS(130), OKO=>SUB_OKOS(130), D=>SUB_DS(130), SO=>SUB_SOS(130));
	DIV131: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(98), SI=>SUB_SOS(99), BI=>SUB_BOS(130), OKI=>SUB_OKOS(132), BO=>SUB_BOS(131), OKO=>SUB_OKOS(131), D=>SUB_DS(131), SO=>SUB_SOS(131));
	DIV132: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(99), SI=>SUB_SOS(100), BI=>SUB_BOS(131), OKI=>SUB_OKOS(133), BO=>SUB_BOS(132), OKO=>SUB_OKOS(132), D=>SUB_DS(132), SO=>SUB_SOS(132));
	DIV133: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(100), SI=>SUB_SOS(101), BI=>SUB_BOS(132), OKI=>SUB_OKOS(134), BO=>SUB_BOS(133), OKO=>SUB_OKOS(133), D=>SUB_DS(133), SO=>SUB_SOS(133));
	DIV134: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(101), SI=>SUB_SOS(102), BI=>SUB_BOS(133), OKI=>SUB_OKOS(135), BO=>SUB_BOS(134), OKO=>SUB_OKOS(134), D=>SUB_DS(134), SO=>SUB_SOS(134));
	DIV135: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(102), SI=>SUB_SOS(103), BI=>SUB_BOS(134), OKI=>SUB_OKOS(136), BO=>SUB_BOS(135), OKO=>SUB_OKOS(135), D=>SUB_DS(135), SO=>SUB_SOS(135));
	DIV136: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(103), SI=>SUB_SOS(104), BI=>SUB_BOS(135), OKI=>SUB_OKOS(137), BO=>SUB_BOS(136), OKO=>SUB_OKOS(136), D=>SUB_DS(136), SO=>SUB_SOS(136));
	DIV137: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(104), SI=>SUB_SOS(105), BI=>SUB_BOS(136), OKI=>SUB_OKOS(138), BO=>SUB_BOS(137), OKO=>SUB_OKOS(137), D=>SUB_DS(137), SO=>SUB_SOS(137));
	DIV138: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(105), SI=>SUB_SOS(106), BI=>SUB_BOS(137), OKI=>SUB_OKOS(139), BO=>SUB_BOS(138), OKO=>SUB_OKOS(138), D=>SUB_DS(138), SO=>SUB_SOS(138));
	DIV139: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(106), SI=>SUB_SOS(107), BI=>SUB_BOS(138), OKI=>SUB_OKOS(140), BO=>SUB_BOS(139), OKO=>SUB_OKOS(139), D=>SUB_DS(139), SO=>SUB_SOS(139));
	DIV140: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(107), SI=>SUB_SOS(108), BI=>SUB_BOS(139), OKI=>SUB_OKOS(141), BO=>SUB_BOS(140), OKO=>SUB_OKOS(140), D=>SUB_DS(140), SO=>SUB_SOS(140));
	DIV141: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(108), SI=>SUB_SOS(109), BI=>SUB_BOS(140), OKI=>SUB_OKOS(142), BO=>SUB_BOS(141), OKO=>SUB_OKOS(141), D=>SUB_DS(141), SO=>SUB_SOS(141));
	DIV142: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(109), SI=>SUB_SOS(110), BI=>SUB_BOS(141), OKI=>SUB_OKOS(143), BO=>SUB_BOS(142), OKO=>SUB_OKOS(142), D=>SUB_DS(142), SO=>SUB_SOS(142));
	DIV143: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(110), SI=>SUB_SOS(111), BI=>SUB_BOS(142), OKI=>SUB_OKOS(144), BO=>SUB_BOS(143), OKO=>SUB_OKOS(143), D=>SUB_DS(143), SO=>SUB_SOS(143));
	DIV144: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(111), SI=>SUB_SOS(112), BI=>SUB_BOS(143), OKI=>SUB_OKOS(145), BO=>SUB_BOS(144), OKO=>SUB_OKOS(144), D=>SUB_DS(144), SO=>SUB_SOS(144));
	DIV145: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(112), SI=>SUB_SOS(113), BI=>SUB_BOS(144), OKI=>SUB_OKOS(146), BO=>SUB_BOS(145), OKO=>SUB_OKOS(145), D=>SUB_DS(145), SO=>SUB_SOS(145));
	DIV146: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(113), SI=>SUB_SOS(114), BI=>SUB_BOS(145), OKI=>SUB_OKOS(147), BO=>SUB_BOS(146), OKO=>SUB_OKOS(146), D=>SUB_DS(146), SO=>SUB_SOS(146));
	DIV147: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(114), SI=>SUB_SOS(115), BI=>SUB_BOS(146), OKI=>SUB_OKOS(148), BO=>SUB_BOS(147), OKO=>SUB_OKOS(147), D=>SUB_DS(147), SO=>SUB_SOS(147));
	DIV148: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(115), SI=>SUB_SOS(116), BI=>SUB_BOS(147), OKI=>SUB_OKOS(149), BO=>SUB_BOS(148), OKO=>SUB_OKOS(148), D=>SUB_DS(148), SO=>SUB_SOS(148));
	DIV149: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(116), SI=>SUB_SOS(117), BI=>SUB_BOS(148), OKI=>SUB_OKOS(150), BO=>SUB_BOS(149), OKO=>SUB_OKOS(149), D=>SUB_DS(149), SO=>SUB_SOS(149));
	DIV150: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(117), SI=>SUB_SOS(118), BI=>SUB_BOS(149), OKI=>SUB_OKOS(151), BO=>SUB_BOS(150), OKO=>SUB_OKOS(150), D=>SUB_DS(150), SO=>SUB_SOS(150));
	DIV151: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(118), SI=>SUB_SOS(119), BI=>SUB_BOS(150), OKI=>SUB_OKOS(152), BO=>SUB_BOS(151), OKO=>SUB_OKOS(151), D=>SUB_DS(151), SO=>SUB_SOS(151));
	DIV152: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(119), SI=>SUB_SOS(120), BI=>SUB_BOS(151), OKI=>SUB_OKOS(153), BO=>SUB_BOS(152), OKO=>SUB_OKOS(152), D=>SUB_DS(152), SO=>SUB_SOS(152));
	DIV153: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(120), SI=>SUB_SOS(121), BI=>SUB_BOS(152), OKI=>SUB_OKOS(154), BO=>SUB_BOS(153), OKO=>SUB_OKOS(153), D=>SUB_DS(153), SO=>SUB_SOS(153));
	DIV154: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(121), SI=>SUB_SOS(122), BI=>SUB_BOS(153), OKI=>SUB_OKOS(155), BO=>SUB_BOS(154), OKO=>SUB_OKOS(154), D=>SUB_DS(154), SO=>SUB_SOS(154));
	DIV155: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(122), SI=>SUB_SOS(123), BI=>SUB_BOS(154), OKI=>SUB_OKOS(156), BO=>SUB_BOS(155), OKO=>SUB_OKOS(155), D=>SUB_DS(155), SO=>SUB_SOS(155));
	DIV156: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(123), SI=>SUB_SOS(124), BI=>SUB_BOS(155), OKI=>SUB_OKOS(157), BO=>SUB_BOS(156), OKO=>SUB_OKOS(156), D=>SUB_DS(156), SO=>SUB_SOS(156));
	DIV157: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(124), SI=>SUB_SOS(125), BI=>SUB_BOS(156), OKI=>SUB_OKOS(158), BO=>SUB_BOS(157), OKO=>SUB_OKOS(157), D=>SUB_DS(157), SO=>SUB_SOS(157));
	DIV158: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(125), SI=>SUB_SOS(126), BI=>SUB_BOS(157), OKI=>SUB_OKOS(159), BO=>SUB_BOS(158), OKO=>SUB_OKOS(158), D=>SUB_DS(158), SO=>SUB_SOS(158));
	DIV159: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(126), SI=>SUB_SOS(127), BI=>SUB_BOS(158), OKI=>BONS(4), BO=>SUB_BOS(159), OKO=>SUB_OKOS(159), D=>SUB_DS(159), SO=>SUB_SOS(159));

	DIV160: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(26), SI=>SUB_SOS(128), BI=>'0', OKI=>SUB_OKOS(161), BO=>SUB_BOS(160), OKO=>SUB_OKOS(160), D=>SUB_DS(160), SO=>SUB_SOS(160));
	DIV161: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(128), SI=>SUB_SOS(129), BI=>SUB_BOS(160), OKI=>SUB_OKOS(162), BO=>SUB_BOS(161), OKO=>SUB_OKOS(161), D=>SUB_DS(161), SO=>SUB_SOS(161));
	DIV162: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(129), SI=>SUB_SOS(130), BI=>SUB_BOS(161), OKI=>SUB_OKOS(163), BO=>SUB_BOS(162), OKO=>SUB_OKOS(162), D=>SUB_DS(162), SO=>SUB_SOS(162));
	DIV163: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(130), SI=>SUB_SOS(131), BI=>SUB_BOS(162), OKI=>SUB_OKOS(164), BO=>SUB_BOS(163), OKO=>SUB_OKOS(163), D=>SUB_DS(163), SO=>SUB_SOS(163));
	DIV164: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(131), SI=>SUB_SOS(132), BI=>SUB_BOS(163), OKI=>SUB_OKOS(165), BO=>SUB_BOS(164), OKO=>SUB_OKOS(164), D=>SUB_DS(164), SO=>SUB_SOS(164));
	DIV165: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(132), SI=>SUB_SOS(133), BI=>SUB_BOS(164), OKI=>SUB_OKOS(166), BO=>SUB_BOS(165), OKO=>SUB_OKOS(165), D=>SUB_DS(165), SO=>SUB_SOS(165));
	DIV166: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(133), SI=>SUB_SOS(134), BI=>SUB_BOS(165), OKI=>SUB_OKOS(167), BO=>SUB_BOS(166), OKO=>SUB_OKOS(166), D=>SUB_DS(166), SO=>SUB_SOS(166));
	DIV167: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(134), SI=>SUB_SOS(135), BI=>SUB_BOS(166), OKI=>SUB_OKOS(168), BO=>SUB_BOS(167), OKO=>SUB_OKOS(167), D=>SUB_DS(167), SO=>SUB_SOS(167));
	DIV168: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(135), SI=>SUB_SOS(136), BI=>SUB_BOS(167), OKI=>SUB_OKOS(169), BO=>SUB_BOS(168), OKO=>SUB_OKOS(168), D=>SUB_DS(168), SO=>SUB_SOS(168));
	DIV169: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(136), SI=>SUB_SOS(137), BI=>SUB_BOS(168), OKI=>SUB_OKOS(170), BO=>SUB_BOS(169), OKO=>SUB_OKOS(169), D=>SUB_DS(169), SO=>SUB_SOS(169));
	DIV170: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(137), SI=>SUB_SOS(138), BI=>SUB_BOS(169), OKI=>SUB_OKOS(171), BO=>SUB_BOS(170), OKO=>SUB_OKOS(170), D=>SUB_DS(170), SO=>SUB_SOS(170));
	DIV171: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(138), SI=>SUB_SOS(139), BI=>SUB_BOS(170), OKI=>SUB_OKOS(172), BO=>SUB_BOS(171), OKO=>SUB_OKOS(171), D=>SUB_DS(171), SO=>SUB_SOS(171));
	DIV172: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(139), SI=>SUB_SOS(140), BI=>SUB_BOS(171), OKI=>SUB_OKOS(173), BO=>SUB_BOS(172), OKO=>SUB_OKOS(172), D=>SUB_DS(172), SO=>SUB_SOS(172));
	DIV173: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(140), SI=>SUB_SOS(141), BI=>SUB_BOS(172), OKI=>SUB_OKOS(174), BO=>SUB_BOS(173), OKO=>SUB_OKOS(173), D=>SUB_DS(173), SO=>SUB_SOS(173));
	DIV174: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(141), SI=>SUB_SOS(142), BI=>SUB_BOS(173), OKI=>SUB_OKOS(175), BO=>SUB_BOS(174), OKO=>SUB_OKOS(174), D=>SUB_DS(174), SO=>SUB_SOS(174));
	DIV175: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(142), SI=>SUB_SOS(143), BI=>SUB_BOS(174), OKI=>SUB_OKOS(176), BO=>SUB_BOS(175), OKO=>SUB_OKOS(175), D=>SUB_DS(175), SO=>SUB_SOS(175));
	DIV176: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(143), SI=>SUB_SOS(144), BI=>SUB_BOS(175), OKI=>SUB_OKOS(177), BO=>SUB_BOS(176), OKO=>SUB_OKOS(176), D=>SUB_DS(176), SO=>SUB_SOS(176));
	DIV177: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(144), SI=>SUB_SOS(145), BI=>SUB_BOS(176), OKI=>SUB_OKOS(178), BO=>SUB_BOS(177), OKO=>SUB_OKOS(177), D=>SUB_DS(177), SO=>SUB_SOS(177));
	DIV178: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(145), SI=>SUB_SOS(146), BI=>SUB_BOS(177), OKI=>SUB_OKOS(179), BO=>SUB_BOS(178), OKO=>SUB_OKOS(178), D=>SUB_DS(178), SO=>SUB_SOS(178));
	DIV179: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(146), SI=>SUB_SOS(147), BI=>SUB_BOS(178), OKI=>SUB_OKOS(180), BO=>SUB_BOS(179), OKO=>SUB_OKOS(179), D=>SUB_DS(179), SO=>SUB_SOS(179));
	DIV180: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(147), SI=>SUB_SOS(148), BI=>SUB_BOS(179), OKI=>SUB_OKOS(181), BO=>SUB_BOS(180), OKO=>SUB_OKOS(180), D=>SUB_DS(180), SO=>SUB_SOS(180));
	DIV181: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(148), SI=>SUB_SOS(149), BI=>SUB_BOS(180), OKI=>SUB_OKOS(182), BO=>SUB_BOS(181), OKO=>SUB_OKOS(181), D=>SUB_DS(181), SO=>SUB_SOS(181));
	DIV182: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(149), SI=>SUB_SOS(150), BI=>SUB_BOS(181), OKI=>SUB_OKOS(183), BO=>SUB_BOS(182), OKO=>SUB_OKOS(182), D=>SUB_DS(182), SO=>SUB_SOS(182));
	DIV183: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(150), SI=>SUB_SOS(151), BI=>SUB_BOS(182), OKI=>SUB_OKOS(184), BO=>SUB_BOS(183), OKO=>SUB_OKOS(183), D=>SUB_DS(183), SO=>SUB_SOS(183));
	DIV184: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(151), SI=>SUB_SOS(152), BI=>SUB_BOS(183), OKI=>SUB_OKOS(185), BO=>SUB_BOS(184), OKO=>SUB_OKOS(184), D=>SUB_DS(184), SO=>SUB_SOS(184));
	DIV185: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(152), SI=>SUB_SOS(153), BI=>SUB_BOS(184), OKI=>SUB_OKOS(186), BO=>SUB_BOS(185), OKO=>SUB_OKOS(185), D=>SUB_DS(185), SO=>SUB_SOS(185));
	DIV186: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(153), SI=>SUB_SOS(154), BI=>SUB_BOS(185), OKI=>SUB_OKOS(187), BO=>SUB_BOS(186), OKO=>SUB_OKOS(186), D=>SUB_DS(186), SO=>SUB_SOS(186));
	DIV187: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(154), SI=>SUB_SOS(155), BI=>SUB_BOS(186), OKI=>SUB_OKOS(188), BO=>SUB_BOS(187), OKO=>SUB_OKOS(187), D=>SUB_DS(187), SO=>SUB_SOS(187));
	DIV188: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(155), SI=>SUB_SOS(156), BI=>SUB_BOS(187), OKI=>SUB_OKOS(189), BO=>SUB_BOS(188), OKO=>SUB_OKOS(188), D=>SUB_DS(188), SO=>SUB_SOS(188));
	DIV189: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(156), SI=>SUB_SOS(157), BI=>SUB_BOS(188), OKI=>SUB_OKOS(190), BO=>SUB_BOS(189), OKO=>SUB_OKOS(189), D=>SUB_DS(189), SO=>SUB_SOS(189));
	DIV190: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(157), SI=>SUB_SOS(158), BI=>SUB_BOS(189), OKI=>SUB_OKOS(191), BO=>SUB_BOS(190), OKO=>SUB_OKOS(190), D=>SUB_DS(190), SO=>SUB_SOS(190));
	DIV191: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(158), SI=>SUB_SOS(159), BI=>SUB_BOS(190), OKI=>BONS(5), BO=>SUB_BOS(191), OKO=>SUB_OKOS(191), D=>SUB_DS(191), SO=>SUB_SOS(191));

	DIV192: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(25), SI=>SUB_SOS(160), BI=>'0', OKI=>SUB_OKOS(193), BO=>SUB_BOS(192), OKO=>SUB_OKOS(192), D=>SUB_DS(192), SO=>SUB_SOS(192));
	DIV193: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(160), SI=>SUB_SOS(161), BI=>SUB_BOS(192), OKI=>SUB_OKOS(194), BO=>SUB_BOS(193), OKO=>SUB_OKOS(193), D=>SUB_DS(193), SO=>SUB_SOS(193));
	DIV194: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(161), SI=>SUB_SOS(162), BI=>SUB_BOS(193), OKI=>SUB_OKOS(195), BO=>SUB_BOS(194), OKO=>SUB_OKOS(194), D=>SUB_DS(194), SO=>SUB_SOS(194));
	DIV195: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(162), SI=>SUB_SOS(163), BI=>SUB_BOS(194), OKI=>SUB_OKOS(196), BO=>SUB_BOS(195), OKO=>SUB_OKOS(195), D=>SUB_DS(195), SO=>SUB_SOS(195));
	DIV196: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(163), SI=>SUB_SOS(164), BI=>SUB_BOS(195), OKI=>SUB_OKOS(197), BO=>SUB_BOS(196), OKO=>SUB_OKOS(196), D=>SUB_DS(196), SO=>SUB_SOS(196));
	DIV197: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(164), SI=>SUB_SOS(165), BI=>SUB_BOS(196), OKI=>SUB_OKOS(198), BO=>SUB_BOS(197), OKO=>SUB_OKOS(197), D=>SUB_DS(197), SO=>SUB_SOS(197));
	DIV198: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(165), SI=>SUB_SOS(166), BI=>SUB_BOS(197), OKI=>SUB_OKOS(199), BO=>SUB_BOS(198), OKO=>SUB_OKOS(198), D=>SUB_DS(198), SO=>SUB_SOS(198));
	DIV199: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(166), SI=>SUB_SOS(167), BI=>SUB_BOS(198), OKI=>SUB_OKOS(200), BO=>SUB_BOS(199), OKO=>SUB_OKOS(199), D=>SUB_DS(199), SO=>SUB_SOS(199));
	DIV200: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(167), SI=>SUB_SOS(168), BI=>SUB_BOS(199), OKI=>SUB_OKOS(201), BO=>SUB_BOS(200), OKO=>SUB_OKOS(200), D=>SUB_DS(200), SO=>SUB_SOS(200));
	DIV201: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(168), SI=>SUB_SOS(169), BI=>SUB_BOS(200), OKI=>SUB_OKOS(202), BO=>SUB_BOS(201), OKO=>SUB_OKOS(201), D=>SUB_DS(201), SO=>SUB_SOS(201));
	DIV202: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(169), SI=>SUB_SOS(170), BI=>SUB_BOS(201), OKI=>SUB_OKOS(203), BO=>SUB_BOS(202), OKO=>SUB_OKOS(202), D=>SUB_DS(202), SO=>SUB_SOS(202));
	DIV203: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(170), SI=>SUB_SOS(171), BI=>SUB_BOS(202), OKI=>SUB_OKOS(204), BO=>SUB_BOS(203), OKO=>SUB_OKOS(203), D=>SUB_DS(203), SO=>SUB_SOS(203));
	DIV204: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(171), SI=>SUB_SOS(172), BI=>SUB_BOS(203), OKI=>SUB_OKOS(205), BO=>SUB_BOS(204), OKO=>SUB_OKOS(204), D=>SUB_DS(204), SO=>SUB_SOS(204));
	DIV205: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(172), SI=>SUB_SOS(173), BI=>SUB_BOS(204), OKI=>SUB_OKOS(206), BO=>SUB_BOS(205), OKO=>SUB_OKOS(205), D=>SUB_DS(205), SO=>SUB_SOS(205));
	DIV206: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(173), SI=>SUB_SOS(174), BI=>SUB_BOS(205), OKI=>SUB_OKOS(207), BO=>SUB_BOS(206), OKO=>SUB_OKOS(206), D=>SUB_DS(206), SO=>SUB_SOS(206));
	DIV207: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(174), SI=>SUB_SOS(175), BI=>SUB_BOS(206), OKI=>SUB_OKOS(208), BO=>SUB_BOS(207), OKO=>SUB_OKOS(207), D=>SUB_DS(207), SO=>SUB_SOS(207));
	DIV208: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(175), SI=>SUB_SOS(176), BI=>SUB_BOS(207), OKI=>SUB_OKOS(209), BO=>SUB_BOS(208), OKO=>SUB_OKOS(208), D=>SUB_DS(208), SO=>SUB_SOS(208));
	DIV209: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(176), SI=>SUB_SOS(177), BI=>SUB_BOS(208), OKI=>SUB_OKOS(210), BO=>SUB_BOS(209), OKO=>SUB_OKOS(209), D=>SUB_DS(209), SO=>SUB_SOS(209));
	DIV210: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(177), SI=>SUB_SOS(178), BI=>SUB_BOS(209), OKI=>SUB_OKOS(211), BO=>SUB_BOS(210), OKO=>SUB_OKOS(210), D=>SUB_DS(210), SO=>SUB_SOS(210));
	DIV211: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(178), SI=>SUB_SOS(179), BI=>SUB_BOS(210), OKI=>SUB_OKOS(212), BO=>SUB_BOS(211), OKO=>SUB_OKOS(211), D=>SUB_DS(211), SO=>SUB_SOS(211));
	DIV212: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(179), SI=>SUB_SOS(180), BI=>SUB_BOS(211), OKI=>SUB_OKOS(213), BO=>SUB_BOS(212), OKO=>SUB_OKOS(212), D=>SUB_DS(212), SO=>SUB_SOS(212));
	DIV213: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(180), SI=>SUB_SOS(181), BI=>SUB_BOS(212), OKI=>SUB_OKOS(214), BO=>SUB_BOS(213), OKO=>SUB_OKOS(213), D=>SUB_DS(213), SO=>SUB_SOS(213));
	DIV214: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(181), SI=>SUB_SOS(182), BI=>SUB_BOS(213), OKI=>SUB_OKOS(215), BO=>SUB_BOS(214), OKO=>SUB_OKOS(214), D=>SUB_DS(214), SO=>SUB_SOS(214));
	DIV215: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(182), SI=>SUB_SOS(183), BI=>SUB_BOS(214), OKI=>SUB_OKOS(216), BO=>SUB_BOS(215), OKO=>SUB_OKOS(215), D=>SUB_DS(215), SO=>SUB_SOS(215));
	DIV216: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(183), SI=>SUB_SOS(184), BI=>SUB_BOS(215), OKI=>SUB_OKOS(217), BO=>SUB_BOS(216), OKO=>SUB_OKOS(216), D=>SUB_DS(216), SO=>SUB_SOS(216));
	DIV217: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(184), SI=>SUB_SOS(185), BI=>SUB_BOS(216), OKI=>SUB_OKOS(218), BO=>SUB_BOS(217), OKO=>SUB_OKOS(217), D=>SUB_DS(217), SO=>SUB_SOS(217));
	DIV218: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(185), SI=>SUB_SOS(186), BI=>SUB_BOS(217), OKI=>SUB_OKOS(219), BO=>SUB_BOS(218), OKO=>SUB_OKOS(218), D=>SUB_DS(218), SO=>SUB_SOS(218));
	DIV219: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(186), SI=>SUB_SOS(187), BI=>SUB_BOS(218), OKI=>SUB_OKOS(220), BO=>SUB_BOS(219), OKO=>SUB_OKOS(219), D=>SUB_DS(219), SO=>SUB_SOS(219));
	DIV220: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(187), SI=>SUB_SOS(188), BI=>SUB_BOS(219), OKI=>SUB_OKOS(221), BO=>SUB_BOS(220), OKO=>SUB_OKOS(220), D=>SUB_DS(220), SO=>SUB_SOS(220));
	DIV221: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(188), SI=>SUB_SOS(189), BI=>SUB_BOS(220), OKI=>SUB_OKOS(222), BO=>SUB_BOS(221), OKO=>SUB_OKOS(221), D=>SUB_DS(221), SO=>SUB_SOS(221));
	DIV222: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(189), SI=>SUB_SOS(190), BI=>SUB_BOS(221), OKI=>SUB_OKOS(223), BO=>SUB_BOS(222), OKO=>SUB_OKOS(222), D=>SUB_DS(222), SO=>SUB_SOS(222));
	DIV223: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(190), SI=>SUB_SOS(191), BI=>SUB_BOS(222), OKI=>BONS(6), BO=>SUB_BOS(223), OKO=>SUB_OKOS(223), D=>SUB_DS(223), SO=>SUB_SOS(223));

	DIV224: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(24), SI=>SUB_SOS(192), BI=>'0', OKI=>SUB_OKOS(225), BO=>SUB_BOS(224), OKO=>SUB_OKOS(224), D=>SUB_DS(224), SO=>SUB_SOS(224));
	DIV225: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(192), SI=>SUB_SOS(193), BI=>SUB_BOS(224), OKI=>SUB_OKOS(226), BO=>SUB_BOS(225), OKO=>SUB_OKOS(225), D=>SUB_DS(225), SO=>SUB_SOS(225));
	DIV226: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(193), SI=>SUB_SOS(194), BI=>SUB_BOS(225), OKI=>SUB_OKOS(227), BO=>SUB_BOS(226), OKO=>SUB_OKOS(226), D=>SUB_DS(226), SO=>SUB_SOS(226));
	DIV227: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(194), SI=>SUB_SOS(195), BI=>SUB_BOS(226), OKI=>SUB_OKOS(228), BO=>SUB_BOS(227), OKO=>SUB_OKOS(227), D=>SUB_DS(227), SO=>SUB_SOS(227));
	DIV228: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(195), SI=>SUB_SOS(196), BI=>SUB_BOS(227), OKI=>SUB_OKOS(229), BO=>SUB_BOS(228), OKO=>SUB_OKOS(228), D=>SUB_DS(228), SO=>SUB_SOS(228));
	DIV229: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(196), SI=>SUB_SOS(197), BI=>SUB_BOS(228), OKI=>SUB_OKOS(230), BO=>SUB_BOS(229), OKO=>SUB_OKOS(229), D=>SUB_DS(229), SO=>SUB_SOS(229));
	DIV230: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(197), SI=>SUB_SOS(198), BI=>SUB_BOS(229), OKI=>SUB_OKOS(231), BO=>SUB_BOS(230), OKO=>SUB_OKOS(230), D=>SUB_DS(230), SO=>SUB_SOS(230));
	DIV231: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(198), SI=>SUB_SOS(199), BI=>SUB_BOS(230), OKI=>SUB_OKOS(232), BO=>SUB_BOS(231), OKO=>SUB_OKOS(231), D=>SUB_DS(231), SO=>SUB_SOS(231));
	DIV232: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(199), SI=>SUB_SOS(200), BI=>SUB_BOS(231), OKI=>SUB_OKOS(233), BO=>SUB_BOS(232), OKO=>SUB_OKOS(232), D=>SUB_DS(232), SO=>SUB_SOS(232));
	DIV233: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(200), SI=>SUB_SOS(201), BI=>SUB_BOS(232), OKI=>SUB_OKOS(234), BO=>SUB_BOS(233), OKO=>SUB_OKOS(233), D=>SUB_DS(233), SO=>SUB_SOS(233));
	DIV234: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(201), SI=>SUB_SOS(202), BI=>SUB_BOS(233), OKI=>SUB_OKOS(235), BO=>SUB_BOS(234), OKO=>SUB_OKOS(234), D=>SUB_DS(234), SO=>SUB_SOS(234));
	DIV235: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(202), SI=>SUB_SOS(203), BI=>SUB_BOS(234), OKI=>SUB_OKOS(236), BO=>SUB_BOS(235), OKO=>SUB_OKOS(235), D=>SUB_DS(235), SO=>SUB_SOS(235));
	DIV236: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(203), SI=>SUB_SOS(204), BI=>SUB_BOS(235), OKI=>SUB_OKOS(237), BO=>SUB_BOS(236), OKO=>SUB_OKOS(236), D=>SUB_DS(236), SO=>SUB_SOS(236));
	DIV237: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(204), SI=>SUB_SOS(205), BI=>SUB_BOS(236), OKI=>SUB_OKOS(238), BO=>SUB_BOS(237), OKO=>SUB_OKOS(237), D=>SUB_DS(237), SO=>SUB_SOS(237));
	DIV238: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(205), SI=>SUB_SOS(206), BI=>SUB_BOS(237), OKI=>SUB_OKOS(239), BO=>SUB_BOS(238), OKO=>SUB_OKOS(238), D=>SUB_DS(238), SO=>SUB_SOS(238));
	DIV239: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(206), SI=>SUB_SOS(207), BI=>SUB_BOS(238), OKI=>SUB_OKOS(240), BO=>SUB_BOS(239), OKO=>SUB_OKOS(239), D=>SUB_DS(239), SO=>SUB_SOS(239));
	DIV240: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(207), SI=>SUB_SOS(208), BI=>SUB_BOS(239), OKI=>SUB_OKOS(241), BO=>SUB_BOS(240), OKO=>SUB_OKOS(240), D=>SUB_DS(240), SO=>SUB_SOS(240));
	DIV241: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(208), SI=>SUB_SOS(209), BI=>SUB_BOS(240), OKI=>SUB_OKOS(242), BO=>SUB_BOS(241), OKO=>SUB_OKOS(241), D=>SUB_DS(241), SO=>SUB_SOS(241));
	DIV242: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(209), SI=>SUB_SOS(210), BI=>SUB_BOS(241), OKI=>SUB_OKOS(243), BO=>SUB_BOS(242), OKO=>SUB_OKOS(242), D=>SUB_DS(242), SO=>SUB_SOS(242));
	DIV243: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(210), SI=>SUB_SOS(211), BI=>SUB_BOS(242), OKI=>SUB_OKOS(244), BO=>SUB_BOS(243), OKO=>SUB_OKOS(243), D=>SUB_DS(243), SO=>SUB_SOS(243));
	DIV244: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(211), SI=>SUB_SOS(212), BI=>SUB_BOS(243), OKI=>SUB_OKOS(245), BO=>SUB_BOS(244), OKO=>SUB_OKOS(244), D=>SUB_DS(244), SO=>SUB_SOS(244));
	DIV245: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(212), SI=>SUB_SOS(213), BI=>SUB_BOS(244), OKI=>SUB_OKOS(246), BO=>SUB_BOS(245), OKO=>SUB_OKOS(245), D=>SUB_DS(245), SO=>SUB_SOS(245));
	DIV246: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(213), SI=>SUB_SOS(214), BI=>SUB_BOS(245), OKI=>SUB_OKOS(247), BO=>SUB_BOS(246), OKO=>SUB_OKOS(246), D=>SUB_DS(246), SO=>SUB_SOS(246));
	DIV247: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(214), SI=>SUB_SOS(215), BI=>SUB_BOS(246), OKI=>SUB_OKOS(248), BO=>SUB_BOS(247), OKO=>SUB_OKOS(247), D=>SUB_DS(247), SO=>SUB_SOS(247));
	DIV248: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(215), SI=>SUB_SOS(216), BI=>SUB_BOS(247), OKI=>SUB_OKOS(249), BO=>SUB_BOS(248), OKO=>SUB_OKOS(248), D=>SUB_DS(248), SO=>SUB_SOS(248));
	DIV249: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(216), SI=>SUB_SOS(217), BI=>SUB_BOS(248), OKI=>SUB_OKOS(250), BO=>SUB_BOS(249), OKO=>SUB_OKOS(249), D=>SUB_DS(249), SO=>SUB_SOS(249));
	DIV250: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(217), SI=>SUB_SOS(218), BI=>SUB_BOS(249), OKI=>SUB_OKOS(251), BO=>SUB_BOS(250), OKO=>SUB_OKOS(250), D=>SUB_DS(250), SO=>SUB_SOS(250));
	DIV251: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(218), SI=>SUB_SOS(219), BI=>SUB_BOS(250), OKI=>SUB_OKOS(252), BO=>SUB_BOS(251), OKO=>SUB_OKOS(251), D=>SUB_DS(251), SO=>SUB_SOS(251));
	DIV252: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(219), SI=>SUB_SOS(220), BI=>SUB_BOS(251), OKI=>SUB_OKOS(253), BO=>SUB_BOS(252), OKO=>SUB_OKOS(252), D=>SUB_DS(252), SO=>SUB_SOS(252));
	DIV253: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(220), SI=>SUB_SOS(221), BI=>SUB_BOS(252), OKI=>SUB_OKOS(254), BO=>SUB_BOS(253), OKO=>SUB_OKOS(253), D=>SUB_DS(253), SO=>SUB_SOS(253));
	DIV254: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(221), SI=>SUB_SOS(222), BI=>SUB_BOS(253), OKI=>SUB_OKOS(255), BO=>SUB_BOS(254), OKO=>SUB_OKOS(254), D=>SUB_DS(254), SO=>SUB_SOS(254));
	DIV255: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(222), SI=>SUB_SOS(223), BI=>SUB_BOS(254), OKI=>BONS(7), BO=>SUB_BOS(255), OKO=>SUB_OKOS(255), D=>SUB_DS(255), SO=>SUB_SOS(255));

	DIV256: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(23), SI=>SUB_SOS(224), BI=>'0', OKI=>SUB_OKOS(257), BO=>SUB_BOS(256), OKO=>SUB_OKOS(256), D=>SUB_DS(256), SO=>SUB_SOS(256));
	DIV257: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(224), SI=>SUB_SOS(225), BI=>SUB_BOS(256), OKI=>SUB_OKOS(258), BO=>SUB_BOS(257), OKO=>SUB_OKOS(257), D=>SUB_DS(257), SO=>SUB_SOS(257));
	DIV258: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(225), SI=>SUB_SOS(226), BI=>SUB_BOS(257), OKI=>SUB_OKOS(259), BO=>SUB_BOS(258), OKO=>SUB_OKOS(258), D=>SUB_DS(258), SO=>SUB_SOS(258));
	DIV259: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(226), SI=>SUB_SOS(227), BI=>SUB_BOS(258), OKI=>SUB_OKOS(260), BO=>SUB_BOS(259), OKO=>SUB_OKOS(259), D=>SUB_DS(259), SO=>SUB_SOS(259));
	DIV260: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(227), SI=>SUB_SOS(228), BI=>SUB_BOS(259), OKI=>SUB_OKOS(261), BO=>SUB_BOS(260), OKO=>SUB_OKOS(260), D=>SUB_DS(260), SO=>SUB_SOS(260));
	DIV261: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(228), SI=>SUB_SOS(229), BI=>SUB_BOS(260), OKI=>SUB_OKOS(262), BO=>SUB_BOS(261), OKO=>SUB_OKOS(261), D=>SUB_DS(261), SO=>SUB_SOS(261));
	DIV262: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(229), SI=>SUB_SOS(230), BI=>SUB_BOS(261), OKI=>SUB_OKOS(263), BO=>SUB_BOS(262), OKO=>SUB_OKOS(262), D=>SUB_DS(262), SO=>SUB_SOS(262));
	DIV263: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(230), SI=>SUB_SOS(231), BI=>SUB_BOS(262), OKI=>SUB_OKOS(264), BO=>SUB_BOS(263), OKO=>SUB_OKOS(263), D=>SUB_DS(263), SO=>SUB_SOS(263));
	DIV264: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(231), SI=>SUB_SOS(232), BI=>SUB_BOS(263), OKI=>SUB_OKOS(265), BO=>SUB_BOS(264), OKO=>SUB_OKOS(264), D=>SUB_DS(264), SO=>SUB_SOS(264));
	DIV265: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(232), SI=>SUB_SOS(233), BI=>SUB_BOS(264), OKI=>SUB_OKOS(266), BO=>SUB_BOS(265), OKO=>SUB_OKOS(265), D=>SUB_DS(265), SO=>SUB_SOS(265));
	DIV266: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(233), SI=>SUB_SOS(234), BI=>SUB_BOS(265), OKI=>SUB_OKOS(267), BO=>SUB_BOS(266), OKO=>SUB_OKOS(266), D=>SUB_DS(266), SO=>SUB_SOS(266));
	DIV267: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(234), SI=>SUB_SOS(235), BI=>SUB_BOS(266), OKI=>SUB_OKOS(268), BO=>SUB_BOS(267), OKO=>SUB_OKOS(267), D=>SUB_DS(267), SO=>SUB_SOS(267));
	DIV268: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(235), SI=>SUB_SOS(236), BI=>SUB_BOS(267), OKI=>SUB_OKOS(269), BO=>SUB_BOS(268), OKO=>SUB_OKOS(268), D=>SUB_DS(268), SO=>SUB_SOS(268));
	DIV269: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(236), SI=>SUB_SOS(237), BI=>SUB_BOS(268), OKI=>SUB_OKOS(270), BO=>SUB_BOS(269), OKO=>SUB_OKOS(269), D=>SUB_DS(269), SO=>SUB_SOS(269));
	DIV270: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(237), SI=>SUB_SOS(238), BI=>SUB_BOS(269), OKI=>SUB_OKOS(271), BO=>SUB_BOS(270), OKO=>SUB_OKOS(270), D=>SUB_DS(270), SO=>SUB_SOS(270));
	DIV271: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(238), SI=>SUB_SOS(239), BI=>SUB_BOS(270), OKI=>SUB_OKOS(272), BO=>SUB_BOS(271), OKO=>SUB_OKOS(271), D=>SUB_DS(271), SO=>SUB_SOS(271));
	DIV272: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(239), SI=>SUB_SOS(240), BI=>SUB_BOS(271), OKI=>SUB_OKOS(273), BO=>SUB_BOS(272), OKO=>SUB_OKOS(272), D=>SUB_DS(272), SO=>SUB_SOS(272));
	DIV273: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(240), SI=>SUB_SOS(241), BI=>SUB_BOS(272), OKI=>SUB_OKOS(274), BO=>SUB_BOS(273), OKO=>SUB_OKOS(273), D=>SUB_DS(273), SO=>SUB_SOS(273));
	DIV274: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(241), SI=>SUB_SOS(242), BI=>SUB_BOS(273), OKI=>SUB_OKOS(275), BO=>SUB_BOS(274), OKO=>SUB_OKOS(274), D=>SUB_DS(274), SO=>SUB_SOS(274));
	DIV275: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(242), SI=>SUB_SOS(243), BI=>SUB_BOS(274), OKI=>SUB_OKOS(276), BO=>SUB_BOS(275), OKO=>SUB_OKOS(275), D=>SUB_DS(275), SO=>SUB_SOS(275));
	DIV276: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(243), SI=>SUB_SOS(244), BI=>SUB_BOS(275), OKI=>SUB_OKOS(277), BO=>SUB_BOS(276), OKO=>SUB_OKOS(276), D=>SUB_DS(276), SO=>SUB_SOS(276));
	DIV277: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(244), SI=>SUB_SOS(245), BI=>SUB_BOS(276), OKI=>SUB_OKOS(278), BO=>SUB_BOS(277), OKO=>SUB_OKOS(277), D=>SUB_DS(277), SO=>SUB_SOS(277));
	DIV278: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(245), SI=>SUB_SOS(246), BI=>SUB_BOS(277), OKI=>SUB_OKOS(279), BO=>SUB_BOS(278), OKO=>SUB_OKOS(278), D=>SUB_DS(278), SO=>SUB_SOS(278));
	DIV279: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(246), SI=>SUB_SOS(247), BI=>SUB_BOS(278), OKI=>SUB_OKOS(280), BO=>SUB_BOS(279), OKO=>SUB_OKOS(279), D=>SUB_DS(279), SO=>SUB_SOS(279));
	DIV280: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(247), SI=>SUB_SOS(248), BI=>SUB_BOS(279), OKI=>SUB_OKOS(281), BO=>SUB_BOS(280), OKO=>SUB_OKOS(280), D=>SUB_DS(280), SO=>SUB_SOS(280));
	DIV281: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(248), SI=>SUB_SOS(249), BI=>SUB_BOS(280), OKI=>SUB_OKOS(282), BO=>SUB_BOS(281), OKO=>SUB_OKOS(281), D=>SUB_DS(281), SO=>SUB_SOS(281));
	DIV282: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(249), SI=>SUB_SOS(250), BI=>SUB_BOS(281), OKI=>SUB_OKOS(283), BO=>SUB_BOS(282), OKO=>SUB_OKOS(282), D=>SUB_DS(282), SO=>SUB_SOS(282));
	DIV283: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(250), SI=>SUB_SOS(251), BI=>SUB_BOS(282), OKI=>SUB_OKOS(284), BO=>SUB_BOS(283), OKO=>SUB_OKOS(283), D=>SUB_DS(283), SO=>SUB_SOS(283));
	DIV284: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(251), SI=>SUB_SOS(252), BI=>SUB_BOS(283), OKI=>SUB_OKOS(285), BO=>SUB_BOS(284), OKO=>SUB_OKOS(284), D=>SUB_DS(284), SO=>SUB_SOS(284));
	DIV285: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(252), SI=>SUB_SOS(253), BI=>SUB_BOS(284), OKI=>SUB_OKOS(286), BO=>SUB_BOS(285), OKO=>SUB_OKOS(285), D=>SUB_DS(285), SO=>SUB_SOS(285));
	DIV286: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(253), SI=>SUB_SOS(254), BI=>SUB_BOS(285), OKI=>SUB_OKOS(287), BO=>SUB_BOS(286), OKO=>SUB_OKOS(286), D=>SUB_DS(286), SO=>SUB_SOS(286));
	DIV287: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(254), SI=>SUB_SOS(255), BI=>SUB_BOS(286), OKI=>BONS(8), BO=>SUB_BOS(287), OKO=>SUB_OKOS(287), D=>SUB_DS(287), SO=>SUB_SOS(287));

	DIV288: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(22), SI=>SUB_SOS(256), BI=>'0', OKI=>SUB_OKOS(289), BO=>SUB_BOS(288), OKO=>SUB_OKOS(288), D=>SUB_DS(288), SO=>SUB_SOS(288));
	DIV289: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(256), SI=>SUB_SOS(257), BI=>SUB_BOS(288), OKI=>SUB_OKOS(290), BO=>SUB_BOS(289), OKO=>SUB_OKOS(289), D=>SUB_DS(289), SO=>SUB_SOS(289));
	DIV290: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(257), SI=>SUB_SOS(258), BI=>SUB_BOS(289), OKI=>SUB_OKOS(291), BO=>SUB_BOS(290), OKO=>SUB_OKOS(290), D=>SUB_DS(290), SO=>SUB_SOS(290));
	DIV291: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(258), SI=>SUB_SOS(259), BI=>SUB_BOS(290), OKI=>SUB_OKOS(292), BO=>SUB_BOS(291), OKO=>SUB_OKOS(291), D=>SUB_DS(291), SO=>SUB_SOS(291));
	DIV292: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(259), SI=>SUB_SOS(260), BI=>SUB_BOS(291), OKI=>SUB_OKOS(293), BO=>SUB_BOS(292), OKO=>SUB_OKOS(292), D=>SUB_DS(292), SO=>SUB_SOS(292));
	DIV293: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(260), SI=>SUB_SOS(261), BI=>SUB_BOS(292), OKI=>SUB_OKOS(294), BO=>SUB_BOS(293), OKO=>SUB_OKOS(293), D=>SUB_DS(293), SO=>SUB_SOS(293));
	DIV294: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(261), SI=>SUB_SOS(262), BI=>SUB_BOS(293), OKI=>SUB_OKOS(295), BO=>SUB_BOS(294), OKO=>SUB_OKOS(294), D=>SUB_DS(294), SO=>SUB_SOS(294));
	DIV295: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(262), SI=>SUB_SOS(263), BI=>SUB_BOS(294), OKI=>SUB_OKOS(296), BO=>SUB_BOS(295), OKO=>SUB_OKOS(295), D=>SUB_DS(295), SO=>SUB_SOS(295));
	DIV296: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(263), SI=>SUB_SOS(264), BI=>SUB_BOS(295), OKI=>SUB_OKOS(297), BO=>SUB_BOS(296), OKO=>SUB_OKOS(296), D=>SUB_DS(296), SO=>SUB_SOS(296));
	DIV297: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(264), SI=>SUB_SOS(265), BI=>SUB_BOS(296), OKI=>SUB_OKOS(298), BO=>SUB_BOS(297), OKO=>SUB_OKOS(297), D=>SUB_DS(297), SO=>SUB_SOS(297));
	DIV298: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(265), SI=>SUB_SOS(266), BI=>SUB_BOS(297), OKI=>SUB_OKOS(299), BO=>SUB_BOS(298), OKO=>SUB_OKOS(298), D=>SUB_DS(298), SO=>SUB_SOS(298));
	DIV299: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(266), SI=>SUB_SOS(267), BI=>SUB_BOS(298), OKI=>SUB_OKOS(300), BO=>SUB_BOS(299), OKO=>SUB_OKOS(299), D=>SUB_DS(299), SO=>SUB_SOS(299));
	DIV300: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(267), SI=>SUB_SOS(268), BI=>SUB_BOS(299), OKI=>SUB_OKOS(301), BO=>SUB_BOS(300), OKO=>SUB_OKOS(300), D=>SUB_DS(300), SO=>SUB_SOS(300));
	DIV301: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(268), SI=>SUB_SOS(269), BI=>SUB_BOS(300), OKI=>SUB_OKOS(302), BO=>SUB_BOS(301), OKO=>SUB_OKOS(301), D=>SUB_DS(301), SO=>SUB_SOS(301));
	DIV302: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(269), SI=>SUB_SOS(270), BI=>SUB_BOS(301), OKI=>SUB_OKOS(303), BO=>SUB_BOS(302), OKO=>SUB_OKOS(302), D=>SUB_DS(302), SO=>SUB_SOS(302));
	DIV303: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(270), SI=>SUB_SOS(271), BI=>SUB_BOS(302), OKI=>SUB_OKOS(304), BO=>SUB_BOS(303), OKO=>SUB_OKOS(303), D=>SUB_DS(303), SO=>SUB_SOS(303));
	DIV304: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(271), SI=>SUB_SOS(272), BI=>SUB_BOS(303), OKI=>SUB_OKOS(305), BO=>SUB_BOS(304), OKO=>SUB_OKOS(304), D=>SUB_DS(304), SO=>SUB_SOS(304));
	DIV305: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(272), SI=>SUB_SOS(273), BI=>SUB_BOS(304), OKI=>SUB_OKOS(306), BO=>SUB_BOS(305), OKO=>SUB_OKOS(305), D=>SUB_DS(305), SO=>SUB_SOS(305));
	DIV306: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(273), SI=>SUB_SOS(274), BI=>SUB_BOS(305), OKI=>SUB_OKOS(307), BO=>SUB_BOS(306), OKO=>SUB_OKOS(306), D=>SUB_DS(306), SO=>SUB_SOS(306));
	DIV307: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(274), SI=>SUB_SOS(275), BI=>SUB_BOS(306), OKI=>SUB_OKOS(308), BO=>SUB_BOS(307), OKO=>SUB_OKOS(307), D=>SUB_DS(307), SO=>SUB_SOS(307));
	DIV308: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(275), SI=>SUB_SOS(276), BI=>SUB_BOS(307), OKI=>SUB_OKOS(309), BO=>SUB_BOS(308), OKO=>SUB_OKOS(308), D=>SUB_DS(308), SO=>SUB_SOS(308));
	DIV309: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(276), SI=>SUB_SOS(277), BI=>SUB_BOS(308), OKI=>SUB_OKOS(310), BO=>SUB_BOS(309), OKO=>SUB_OKOS(309), D=>SUB_DS(309), SO=>SUB_SOS(309));
	DIV310: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(277), SI=>SUB_SOS(278), BI=>SUB_BOS(309), OKI=>SUB_OKOS(311), BO=>SUB_BOS(310), OKO=>SUB_OKOS(310), D=>SUB_DS(310), SO=>SUB_SOS(310));
	DIV311: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(278), SI=>SUB_SOS(279), BI=>SUB_BOS(310), OKI=>SUB_OKOS(312), BO=>SUB_BOS(311), OKO=>SUB_OKOS(311), D=>SUB_DS(311), SO=>SUB_SOS(311));
	DIV312: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(279), SI=>SUB_SOS(280), BI=>SUB_BOS(311), OKI=>SUB_OKOS(313), BO=>SUB_BOS(312), OKO=>SUB_OKOS(312), D=>SUB_DS(312), SO=>SUB_SOS(312));
	DIV313: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(280), SI=>SUB_SOS(281), BI=>SUB_BOS(312), OKI=>SUB_OKOS(314), BO=>SUB_BOS(313), OKO=>SUB_OKOS(313), D=>SUB_DS(313), SO=>SUB_SOS(313));
	DIV314: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(281), SI=>SUB_SOS(282), BI=>SUB_BOS(313), OKI=>SUB_OKOS(315), BO=>SUB_BOS(314), OKO=>SUB_OKOS(314), D=>SUB_DS(314), SO=>SUB_SOS(314));
	DIV315: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(282), SI=>SUB_SOS(283), BI=>SUB_BOS(314), OKI=>SUB_OKOS(316), BO=>SUB_BOS(315), OKO=>SUB_OKOS(315), D=>SUB_DS(315), SO=>SUB_SOS(315));
	DIV316: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(283), SI=>SUB_SOS(284), BI=>SUB_BOS(315), OKI=>SUB_OKOS(317), BO=>SUB_BOS(316), OKO=>SUB_OKOS(316), D=>SUB_DS(316), SO=>SUB_SOS(316));
	DIV317: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(284), SI=>SUB_SOS(285), BI=>SUB_BOS(316), OKI=>SUB_OKOS(318), BO=>SUB_BOS(317), OKO=>SUB_OKOS(317), D=>SUB_DS(317), SO=>SUB_SOS(317));
	DIV318: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(285), SI=>SUB_SOS(286), BI=>SUB_BOS(317), OKI=>SUB_OKOS(319), BO=>SUB_BOS(318), OKO=>SUB_OKOS(318), D=>SUB_DS(318), SO=>SUB_SOS(318));
	DIV319: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(286), SI=>SUB_SOS(287), BI=>SUB_BOS(318), OKI=>BONS(9), BO=>SUB_BOS(319), OKO=>SUB_OKOS(319), D=>SUB_DS(319), SO=>SUB_SOS(319));

	DIV320: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(21), SI=>SUB_SOS(288), BI=>'0', OKI=>SUB_OKOS(321), BO=>SUB_BOS(320), OKO=>SUB_OKOS(320), D=>SUB_DS(320), SO=>SUB_SOS(320));
	DIV321: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(288), SI=>SUB_SOS(289), BI=>SUB_BOS(320), OKI=>SUB_OKOS(322), BO=>SUB_BOS(321), OKO=>SUB_OKOS(321), D=>SUB_DS(321), SO=>SUB_SOS(321));
	DIV322: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(289), SI=>SUB_SOS(290), BI=>SUB_BOS(321), OKI=>SUB_OKOS(323), BO=>SUB_BOS(322), OKO=>SUB_OKOS(322), D=>SUB_DS(322), SO=>SUB_SOS(322));
	DIV323: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(290), SI=>SUB_SOS(291), BI=>SUB_BOS(322), OKI=>SUB_OKOS(324), BO=>SUB_BOS(323), OKO=>SUB_OKOS(323), D=>SUB_DS(323), SO=>SUB_SOS(323));
	DIV324: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(291), SI=>SUB_SOS(292), BI=>SUB_BOS(323), OKI=>SUB_OKOS(325), BO=>SUB_BOS(324), OKO=>SUB_OKOS(324), D=>SUB_DS(324), SO=>SUB_SOS(324));
	DIV325: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(292), SI=>SUB_SOS(293), BI=>SUB_BOS(324), OKI=>SUB_OKOS(326), BO=>SUB_BOS(325), OKO=>SUB_OKOS(325), D=>SUB_DS(325), SO=>SUB_SOS(325));
	DIV326: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(293), SI=>SUB_SOS(294), BI=>SUB_BOS(325), OKI=>SUB_OKOS(327), BO=>SUB_BOS(326), OKO=>SUB_OKOS(326), D=>SUB_DS(326), SO=>SUB_SOS(326));
	DIV327: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(294), SI=>SUB_SOS(295), BI=>SUB_BOS(326), OKI=>SUB_OKOS(328), BO=>SUB_BOS(327), OKO=>SUB_OKOS(327), D=>SUB_DS(327), SO=>SUB_SOS(327));
	DIV328: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(295), SI=>SUB_SOS(296), BI=>SUB_BOS(327), OKI=>SUB_OKOS(329), BO=>SUB_BOS(328), OKO=>SUB_OKOS(328), D=>SUB_DS(328), SO=>SUB_SOS(328));
	DIV329: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(296), SI=>SUB_SOS(297), BI=>SUB_BOS(328), OKI=>SUB_OKOS(330), BO=>SUB_BOS(329), OKO=>SUB_OKOS(329), D=>SUB_DS(329), SO=>SUB_SOS(329));
	DIV330: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(297), SI=>SUB_SOS(298), BI=>SUB_BOS(329), OKI=>SUB_OKOS(331), BO=>SUB_BOS(330), OKO=>SUB_OKOS(330), D=>SUB_DS(330), SO=>SUB_SOS(330));
	DIV331: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(298), SI=>SUB_SOS(299), BI=>SUB_BOS(330), OKI=>SUB_OKOS(332), BO=>SUB_BOS(331), OKO=>SUB_OKOS(331), D=>SUB_DS(331), SO=>SUB_SOS(331));
	DIV332: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(299), SI=>SUB_SOS(300), BI=>SUB_BOS(331), OKI=>SUB_OKOS(333), BO=>SUB_BOS(332), OKO=>SUB_OKOS(332), D=>SUB_DS(332), SO=>SUB_SOS(332));
	DIV333: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(300), SI=>SUB_SOS(301), BI=>SUB_BOS(332), OKI=>SUB_OKOS(334), BO=>SUB_BOS(333), OKO=>SUB_OKOS(333), D=>SUB_DS(333), SO=>SUB_SOS(333));
	DIV334: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(301), SI=>SUB_SOS(302), BI=>SUB_BOS(333), OKI=>SUB_OKOS(335), BO=>SUB_BOS(334), OKO=>SUB_OKOS(334), D=>SUB_DS(334), SO=>SUB_SOS(334));
	DIV335: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(302), SI=>SUB_SOS(303), BI=>SUB_BOS(334), OKI=>SUB_OKOS(336), BO=>SUB_BOS(335), OKO=>SUB_OKOS(335), D=>SUB_DS(335), SO=>SUB_SOS(335));
	DIV336: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(303), SI=>SUB_SOS(304), BI=>SUB_BOS(335), OKI=>SUB_OKOS(337), BO=>SUB_BOS(336), OKO=>SUB_OKOS(336), D=>SUB_DS(336), SO=>SUB_SOS(336));
	DIV337: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(304), SI=>SUB_SOS(305), BI=>SUB_BOS(336), OKI=>SUB_OKOS(338), BO=>SUB_BOS(337), OKO=>SUB_OKOS(337), D=>SUB_DS(337), SO=>SUB_SOS(337));
	DIV338: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(305), SI=>SUB_SOS(306), BI=>SUB_BOS(337), OKI=>SUB_OKOS(339), BO=>SUB_BOS(338), OKO=>SUB_OKOS(338), D=>SUB_DS(338), SO=>SUB_SOS(338));
	DIV339: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(306), SI=>SUB_SOS(307), BI=>SUB_BOS(338), OKI=>SUB_OKOS(340), BO=>SUB_BOS(339), OKO=>SUB_OKOS(339), D=>SUB_DS(339), SO=>SUB_SOS(339));
	DIV340: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(307), SI=>SUB_SOS(308), BI=>SUB_BOS(339), OKI=>SUB_OKOS(341), BO=>SUB_BOS(340), OKO=>SUB_OKOS(340), D=>SUB_DS(340), SO=>SUB_SOS(340));
	DIV341: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(308), SI=>SUB_SOS(309), BI=>SUB_BOS(340), OKI=>SUB_OKOS(342), BO=>SUB_BOS(341), OKO=>SUB_OKOS(341), D=>SUB_DS(341), SO=>SUB_SOS(341));
	DIV342: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(309), SI=>SUB_SOS(310), BI=>SUB_BOS(341), OKI=>SUB_OKOS(343), BO=>SUB_BOS(342), OKO=>SUB_OKOS(342), D=>SUB_DS(342), SO=>SUB_SOS(342));
	DIV343: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(310), SI=>SUB_SOS(311), BI=>SUB_BOS(342), OKI=>SUB_OKOS(344), BO=>SUB_BOS(343), OKO=>SUB_OKOS(343), D=>SUB_DS(343), SO=>SUB_SOS(343));
	DIV344: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(311), SI=>SUB_SOS(312), BI=>SUB_BOS(343), OKI=>SUB_OKOS(345), BO=>SUB_BOS(344), OKO=>SUB_OKOS(344), D=>SUB_DS(344), SO=>SUB_SOS(344));
	DIV345: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(312), SI=>SUB_SOS(313), BI=>SUB_BOS(344), OKI=>SUB_OKOS(346), BO=>SUB_BOS(345), OKO=>SUB_OKOS(345), D=>SUB_DS(345), SO=>SUB_SOS(345));
	DIV346: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(313), SI=>SUB_SOS(314), BI=>SUB_BOS(345), OKI=>SUB_OKOS(347), BO=>SUB_BOS(346), OKO=>SUB_OKOS(346), D=>SUB_DS(346), SO=>SUB_SOS(346));
	DIV347: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(314), SI=>SUB_SOS(315), BI=>SUB_BOS(346), OKI=>SUB_OKOS(348), BO=>SUB_BOS(347), OKO=>SUB_OKOS(347), D=>SUB_DS(347), SO=>SUB_SOS(347));
	DIV348: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(315), SI=>SUB_SOS(316), BI=>SUB_BOS(347), OKI=>SUB_OKOS(349), BO=>SUB_BOS(348), OKO=>SUB_OKOS(348), D=>SUB_DS(348), SO=>SUB_SOS(348));
	DIV349: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(316), SI=>SUB_SOS(317), BI=>SUB_BOS(348), OKI=>SUB_OKOS(350), BO=>SUB_BOS(349), OKO=>SUB_OKOS(349), D=>SUB_DS(349), SO=>SUB_SOS(349));
	DIV350: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(317), SI=>SUB_SOS(318), BI=>SUB_BOS(349), OKI=>SUB_OKOS(351), BO=>SUB_BOS(350), OKO=>SUB_OKOS(350), D=>SUB_DS(350), SO=>SUB_SOS(350));
	DIV351: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(318), SI=>SUB_SOS(319), BI=>SUB_BOS(350), OKI=>BONS(10), BO=>SUB_BOS(351), OKO=>SUB_OKOS(351), D=>SUB_DS(351), SO=>SUB_SOS(351));

	DIV352: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(20), SI=>SUB_SOS(320), BI=>'0', OKI=>SUB_OKOS(353), BO=>SUB_BOS(352), OKO=>SUB_OKOS(352), D=>SUB_DS(352), SO=>SUB_SOS(352));
	DIV353: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(320), SI=>SUB_SOS(321), BI=>SUB_BOS(352), OKI=>SUB_OKOS(354), BO=>SUB_BOS(353), OKO=>SUB_OKOS(353), D=>SUB_DS(353), SO=>SUB_SOS(353));
	DIV354: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(321), SI=>SUB_SOS(322), BI=>SUB_BOS(353), OKI=>SUB_OKOS(355), BO=>SUB_BOS(354), OKO=>SUB_OKOS(354), D=>SUB_DS(354), SO=>SUB_SOS(354));
	DIV355: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(322), SI=>SUB_SOS(323), BI=>SUB_BOS(354), OKI=>SUB_OKOS(356), BO=>SUB_BOS(355), OKO=>SUB_OKOS(355), D=>SUB_DS(355), SO=>SUB_SOS(355));
	DIV356: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(323), SI=>SUB_SOS(324), BI=>SUB_BOS(355), OKI=>SUB_OKOS(357), BO=>SUB_BOS(356), OKO=>SUB_OKOS(356), D=>SUB_DS(356), SO=>SUB_SOS(356));
	DIV357: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(324), SI=>SUB_SOS(325), BI=>SUB_BOS(356), OKI=>SUB_OKOS(358), BO=>SUB_BOS(357), OKO=>SUB_OKOS(357), D=>SUB_DS(357), SO=>SUB_SOS(357));
	DIV358: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(325), SI=>SUB_SOS(326), BI=>SUB_BOS(357), OKI=>SUB_OKOS(359), BO=>SUB_BOS(358), OKO=>SUB_OKOS(358), D=>SUB_DS(358), SO=>SUB_SOS(358));
	DIV359: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(326), SI=>SUB_SOS(327), BI=>SUB_BOS(358), OKI=>SUB_OKOS(360), BO=>SUB_BOS(359), OKO=>SUB_OKOS(359), D=>SUB_DS(359), SO=>SUB_SOS(359));
	DIV360: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(327), SI=>SUB_SOS(328), BI=>SUB_BOS(359), OKI=>SUB_OKOS(361), BO=>SUB_BOS(360), OKO=>SUB_OKOS(360), D=>SUB_DS(360), SO=>SUB_SOS(360));
	DIV361: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(328), SI=>SUB_SOS(329), BI=>SUB_BOS(360), OKI=>SUB_OKOS(362), BO=>SUB_BOS(361), OKO=>SUB_OKOS(361), D=>SUB_DS(361), SO=>SUB_SOS(361));
	DIV362: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(329), SI=>SUB_SOS(330), BI=>SUB_BOS(361), OKI=>SUB_OKOS(363), BO=>SUB_BOS(362), OKO=>SUB_OKOS(362), D=>SUB_DS(362), SO=>SUB_SOS(362));
	DIV363: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(330), SI=>SUB_SOS(331), BI=>SUB_BOS(362), OKI=>SUB_OKOS(364), BO=>SUB_BOS(363), OKO=>SUB_OKOS(363), D=>SUB_DS(363), SO=>SUB_SOS(363));
	DIV364: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(331), SI=>SUB_SOS(332), BI=>SUB_BOS(363), OKI=>SUB_OKOS(365), BO=>SUB_BOS(364), OKO=>SUB_OKOS(364), D=>SUB_DS(364), SO=>SUB_SOS(364));
	DIV365: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(332), SI=>SUB_SOS(333), BI=>SUB_BOS(364), OKI=>SUB_OKOS(366), BO=>SUB_BOS(365), OKO=>SUB_OKOS(365), D=>SUB_DS(365), SO=>SUB_SOS(365));
	DIV366: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(333), SI=>SUB_SOS(334), BI=>SUB_BOS(365), OKI=>SUB_OKOS(367), BO=>SUB_BOS(366), OKO=>SUB_OKOS(366), D=>SUB_DS(366), SO=>SUB_SOS(366));
	DIV367: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(334), SI=>SUB_SOS(335), BI=>SUB_BOS(366), OKI=>SUB_OKOS(368), BO=>SUB_BOS(367), OKO=>SUB_OKOS(367), D=>SUB_DS(367), SO=>SUB_SOS(367));
	DIV368: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(335), SI=>SUB_SOS(336), BI=>SUB_BOS(367), OKI=>SUB_OKOS(369), BO=>SUB_BOS(368), OKO=>SUB_OKOS(368), D=>SUB_DS(368), SO=>SUB_SOS(368));
	DIV369: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(336), SI=>SUB_SOS(337), BI=>SUB_BOS(368), OKI=>SUB_OKOS(370), BO=>SUB_BOS(369), OKO=>SUB_OKOS(369), D=>SUB_DS(369), SO=>SUB_SOS(369));
	DIV370: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(337), SI=>SUB_SOS(338), BI=>SUB_BOS(369), OKI=>SUB_OKOS(371), BO=>SUB_BOS(370), OKO=>SUB_OKOS(370), D=>SUB_DS(370), SO=>SUB_SOS(370));
	DIV371: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(338), SI=>SUB_SOS(339), BI=>SUB_BOS(370), OKI=>SUB_OKOS(372), BO=>SUB_BOS(371), OKO=>SUB_OKOS(371), D=>SUB_DS(371), SO=>SUB_SOS(371));
	DIV372: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(339), SI=>SUB_SOS(340), BI=>SUB_BOS(371), OKI=>SUB_OKOS(373), BO=>SUB_BOS(372), OKO=>SUB_OKOS(372), D=>SUB_DS(372), SO=>SUB_SOS(372));
	DIV373: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(340), SI=>SUB_SOS(341), BI=>SUB_BOS(372), OKI=>SUB_OKOS(374), BO=>SUB_BOS(373), OKO=>SUB_OKOS(373), D=>SUB_DS(373), SO=>SUB_SOS(373));
	DIV374: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(341), SI=>SUB_SOS(342), BI=>SUB_BOS(373), OKI=>SUB_OKOS(375), BO=>SUB_BOS(374), OKO=>SUB_OKOS(374), D=>SUB_DS(374), SO=>SUB_SOS(374));
	DIV375: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(342), SI=>SUB_SOS(343), BI=>SUB_BOS(374), OKI=>SUB_OKOS(376), BO=>SUB_BOS(375), OKO=>SUB_OKOS(375), D=>SUB_DS(375), SO=>SUB_SOS(375));
	DIV376: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(343), SI=>SUB_SOS(344), BI=>SUB_BOS(375), OKI=>SUB_OKOS(377), BO=>SUB_BOS(376), OKO=>SUB_OKOS(376), D=>SUB_DS(376), SO=>SUB_SOS(376));
	DIV377: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(344), SI=>SUB_SOS(345), BI=>SUB_BOS(376), OKI=>SUB_OKOS(378), BO=>SUB_BOS(377), OKO=>SUB_OKOS(377), D=>SUB_DS(377), SO=>SUB_SOS(377));
	DIV378: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(345), SI=>SUB_SOS(346), BI=>SUB_BOS(377), OKI=>SUB_OKOS(379), BO=>SUB_BOS(378), OKO=>SUB_OKOS(378), D=>SUB_DS(378), SO=>SUB_SOS(378));
	DIV379: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(346), SI=>SUB_SOS(347), BI=>SUB_BOS(378), OKI=>SUB_OKOS(380), BO=>SUB_BOS(379), OKO=>SUB_OKOS(379), D=>SUB_DS(379), SO=>SUB_SOS(379));
	DIV380: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(347), SI=>SUB_SOS(348), BI=>SUB_BOS(379), OKI=>SUB_OKOS(381), BO=>SUB_BOS(380), OKO=>SUB_OKOS(380), D=>SUB_DS(380), SO=>SUB_SOS(380));
	DIV381: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(348), SI=>SUB_SOS(349), BI=>SUB_BOS(380), OKI=>SUB_OKOS(382), BO=>SUB_BOS(381), OKO=>SUB_OKOS(381), D=>SUB_DS(381), SO=>SUB_SOS(381));
	DIV382: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(349), SI=>SUB_SOS(350), BI=>SUB_BOS(381), OKI=>SUB_OKOS(383), BO=>SUB_BOS(382), OKO=>SUB_OKOS(382), D=>SUB_DS(382), SO=>SUB_SOS(382));
	DIV383: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(350), SI=>SUB_SOS(351), BI=>SUB_BOS(382), OKI=>BONS(11), BO=>SUB_BOS(383), OKO=>SUB_OKOS(383), D=>SUB_DS(383), SO=>SUB_SOS(383));

	DIV384: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(19), SI=>SUB_SOS(352), BI=>'0', OKI=>SUB_OKOS(385), BO=>SUB_BOS(384), OKO=>SUB_OKOS(384), D=>SUB_DS(384), SO=>SUB_SOS(384));
	DIV385: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(352), SI=>SUB_SOS(353), BI=>SUB_BOS(384), OKI=>SUB_OKOS(386), BO=>SUB_BOS(385), OKO=>SUB_OKOS(385), D=>SUB_DS(385), SO=>SUB_SOS(385));
	DIV386: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(353), SI=>SUB_SOS(354), BI=>SUB_BOS(385), OKI=>SUB_OKOS(387), BO=>SUB_BOS(386), OKO=>SUB_OKOS(386), D=>SUB_DS(386), SO=>SUB_SOS(386));
	DIV387: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(354), SI=>SUB_SOS(355), BI=>SUB_BOS(386), OKI=>SUB_OKOS(388), BO=>SUB_BOS(387), OKO=>SUB_OKOS(387), D=>SUB_DS(387), SO=>SUB_SOS(387));
	DIV388: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(355), SI=>SUB_SOS(356), BI=>SUB_BOS(387), OKI=>SUB_OKOS(389), BO=>SUB_BOS(388), OKO=>SUB_OKOS(388), D=>SUB_DS(388), SO=>SUB_SOS(388));
	DIV389: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(356), SI=>SUB_SOS(357), BI=>SUB_BOS(388), OKI=>SUB_OKOS(390), BO=>SUB_BOS(389), OKO=>SUB_OKOS(389), D=>SUB_DS(389), SO=>SUB_SOS(389));
	DIV390: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(357), SI=>SUB_SOS(358), BI=>SUB_BOS(389), OKI=>SUB_OKOS(391), BO=>SUB_BOS(390), OKO=>SUB_OKOS(390), D=>SUB_DS(390), SO=>SUB_SOS(390));
	DIV391: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(358), SI=>SUB_SOS(359), BI=>SUB_BOS(390), OKI=>SUB_OKOS(392), BO=>SUB_BOS(391), OKO=>SUB_OKOS(391), D=>SUB_DS(391), SO=>SUB_SOS(391));
	DIV392: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(359), SI=>SUB_SOS(360), BI=>SUB_BOS(391), OKI=>SUB_OKOS(393), BO=>SUB_BOS(392), OKO=>SUB_OKOS(392), D=>SUB_DS(392), SO=>SUB_SOS(392));
	DIV393: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(360), SI=>SUB_SOS(361), BI=>SUB_BOS(392), OKI=>SUB_OKOS(394), BO=>SUB_BOS(393), OKO=>SUB_OKOS(393), D=>SUB_DS(393), SO=>SUB_SOS(393));
	DIV394: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(361), SI=>SUB_SOS(362), BI=>SUB_BOS(393), OKI=>SUB_OKOS(395), BO=>SUB_BOS(394), OKO=>SUB_OKOS(394), D=>SUB_DS(394), SO=>SUB_SOS(394));
	DIV395: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(362), SI=>SUB_SOS(363), BI=>SUB_BOS(394), OKI=>SUB_OKOS(396), BO=>SUB_BOS(395), OKO=>SUB_OKOS(395), D=>SUB_DS(395), SO=>SUB_SOS(395));
	DIV396: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(363), SI=>SUB_SOS(364), BI=>SUB_BOS(395), OKI=>SUB_OKOS(397), BO=>SUB_BOS(396), OKO=>SUB_OKOS(396), D=>SUB_DS(396), SO=>SUB_SOS(396));
	DIV397: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(364), SI=>SUB_SOS(365), BI=>SUB_BOS(396), OKI=>SUB_OKOS(398), BO=>SUB_BOS(397), OKO=>SUB_OKOS(397), D=>SUB_DS(397), SO=>SUB_SOS(397));
	DIV398: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(365), SI=>SUB_SOS(366), BI=>SUB_BOS(397), OKI=>SUB_OKOS(399), BO=>SUB_BOS(398), OKO=>SUB_OKOS(398), D=>SUB_DS(398), SO=>SUB_SOS(398));
	DIV399: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(366), SI=>SUB_SOS(367), BI=>SUB_BOS(398), OKI=>SUB_OKOS(400), BO=>SUB_BOS(399), OKO=>SUB_OKOS(399), D=>SUB_DS(399), SO=>SUB_SOS(399));
	DIV400: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(367), SI=>SUB_SOS(368), BI=>SUB_BOS(399), OKI=>SUB_OKOS(401), BO=>SUB_BOS(400), OKO=>SUB_OKOS(400), D=>SUB_DS(400), SO=>SUB_SOS(400));
	DIV401: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(368), SI=>SUB_SOS(369), BI=>SUB_BOS(400), OKI=>SUB_OKOS(402), BO=>SUB_BOS(401), OKO=>SUB_OKOS(401), D=>SUB_DS(401), SO=>SUB_SOS(401));
	DIV402: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(369), SI=>SUB_SOS(370), BI=>SUB_BOS(401), OKI=>SUB_OKOS(403), BO=>SUB_BOS(402), OKO=>SUB_OKOS(402), D=>SUB_DS(402), SO=>SUB_SOS(402));
	DIV403: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(370), SI=>SUB_SOS(371), BI=>SUB_BOS(402), OKI=>SUB_OKOS(404), BO=>SUB_BOS(403), OKO=>SUB_OKOS(403), D=>SUB_DS(403), SO=>SUB_SOS(403));
	DIV404: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(371), SI=>SUB_SOS(372), BI=>SUB_BOS(403), OKI=>SUB_OKOS(405), BO=>SUB_BOS(404), OKO=>SUB_OKOS(404), D=>SUB_DS(404), SO=>SUB_SOS(404));
	DIV405: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(372), SI=>SUB_SOS(373), BI=>SUB_BOS(404), OKI=>SUB_OKOS(406), BO=>SUB_BOS(405), OKO=>SUB_OKOS(405), D=>SUB_DS(405), SO=>SUB_SOS(405));
	DIV406: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(373), SI=>SUB_SOS(374), BI=>SUB_BOS(405), OKI=>SUB_OKOS(407), BO=>SUB_BOS(406), OKO=>SUB_OKOS(406), D=>SUB_DS(406), SO=>SUB_SOS(406));
	DIV407: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(374), SI=>SUB_SOS(375), BI=>SUB_BOS(406), OKI=>SUB_OKOS(408), BO=>SUB_BOS(407), OKO=>SUB_OKOS(407), D=>SUB_DS(407), SO=>SUB_SOS(407));
	DIV408: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(375), SI=>SUB_SOS(376), BI=>SUB_BOS(407), OKI=>SUB_OKOS(409), BO=>SUB_BOS(408), OKO=>SUB_OKOS(408), D=>SUB_DS(408), SO=>SUB_SOS(408));
	DIV409: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(376), SI=>SUB_SOS(377), BI=>SUB_BOS(408), OKI=>SUB_OKOS(410), BO=>SUB_BOS(409), OKO=>SUB_OKOS(409), D=>SUB_DS(409), SO=>SUB_SOS(409));
	DIV410: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(377), SI=>SUB_SOS(378), BI=>SUB_BOS(409), OKI=>SUB_OKOS(411), BO=>SUB_BOS(410), OKO=>SUB_OKOS(410), D=>SUB_DS(410), SO=>SUB_SOS(410));
	DIV411: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(378), SI=>SUB_SOS(379), BI=>SUB_BOS(410), OKI=>SUB_OKOS(412), BO=>SUB_BOS(411), OKO=>SUB_OKOS(411), D=>SUB_DS(411), SO=>SUB_SOS(411));
	DIV412: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(379), SI=>SUB_SOS(380), BI=>SUB_BOS(411), OKI=>SUB_OKOS(413), BO=>SUB_BOS(412), OKO=>SUB_OKOS(412), D=>SUB_DS(412), SO=>SUB_SOS(412));
	DIV413: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(380), SI=>SUB_SOS(381), BI=>SUB_BOS(412), OKI=>SUB_OKOS(414), BO=>SUB_BOS(413), OKO=>SUB_OKOS(413), D=>SUB_DS(413), SO=>SUB_SOS(413));
	DIV414: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(381), SI=>SUB_SOS(382), BI=>SUB_BOS(413), OKI=>SUB_OKOS(415), BO=>SUB_BOS(414), OKO=>SUB_OKOS(414), D=>SUB_DS(414), SO=>SUB_SOS(414));
	DIV415: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(382), SI=>SUB_SOS(383), BI=>SUB_BOS(414), OKI=>BONS(12), BO=>SUB_BOS(415), OKO=>SUB_OKOS(415), D=>SUB_DS(415), SO=>SUB_SOS(415));

	DIV416: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(18), SI=>SUB_SOS(384), BI=>'0', OKI=>SUB_OKOS(417), BO=>SUB_BOS(416), OKO=>SUB_OKOS(416), D=>SUB_DS(416), SO=>SUB_SOS(416));
	DIV417: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(384), SI=>SUB_SOS(385), BI=>SUB_BOS(416), OKI=>SUB_OKOS(418), BO=>SUB_BOS(417), OKO=>SUB_OKOS(417), D=>SUB_DS(417), SO=>SUB_SOS(417));
	DIV418: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(385), SI=>SUB_SOS(386), BI=>SUB_BOS(417), OKI=>SUB_OKOS(419), BO=>SUB_BOS(418), OKO=>SUB_OKOS(418), D=>SUB_DS(418), SO=>SUB_SOS(418));
	DIV419: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(386), SI=>SUB_SOS(387), BI=>SUB_BOS(418), OKI=>SUB_OKOS(420), BO=>SUB_BOS(419), OKO=>SUB_OKOS(419), D=>SUB_DS(419), SO=>SUB_SOS(419));
	DIV420: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(387), SI=>SUB_SOS(388), BI=>SUB_BOS(419), OKI=>SUB_OKOS(421), BO=>SUB_BOS(420), OKO=>SUB_OKOS(420), D=>SUB_DS(420), SO=>SUB_SOS(420));
	DIV421: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(388), SI=>SUB_SOS(389), BI=>SUB_BOS(420), OKI=>SUB_OKOS(422), BO=>SUB_BOS(421), OKO=>SUB_OKOS(421), D=>SUB_DS(421), SO=>SUB_SOS(421));
	DIV422: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(389), SI=>SUB_SOS(390), BI=>SUB_BOS(421), OKI=>SUB_OKOS(423), BO=>SUB_BOS(422), OKO=>SUB_OKOS(422), D=>SUB_DS(422), SO=>SUB_SOS(422));
	DIV423: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(390), SI=>SUB_SOS(391), BI=>SUB_BOS(422), OKI=>SUB_OKOS(424), BO=>SUB_BOS(423), OKO=>SUB_OKOS(423), D=>SUB_DS(423), SO=>SUB_SOS(423));
	DIV424: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(391), SI=>SUB_SOS(392), BI=>SUB_BOS(423), OKI=>SUB_OKOS(425), BO=>SUB_BOS(424), OKO=>SUB_OKOS(424), D=>SUB_DS(424), SO=>SUB_SOS(424));
	DIV425: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(392), SI=>SUB_SOS(393), BI=>SUB_BOS(424), OKI=>SUB_OKOS(426), BO=>SUB_BOS(425), OKO=>SUB_OKOS(425), D=>SUB_DS(425), SO=>SUB_SOS(425));
	DIV426: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(393), SI=>SUB_SOS(394), BI=>SUB_BOS(425), OKI=>SUB_OKOS(427), BO=>SUB_BOS(426), OKO=>SUB_OKOS(426), D=>SUB_DS(426), SO=>SUB_SOS(426));
	DIV427: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(394), SI=>SUB_SOS(395), BI=>SUB_BOS(426), OKI=>SUB_OKOS(428), BO=>SUB_BOS(427), OKO=>SUB_OKOS(427), D=>SUB_DS(427), SO=>SUB_SOS(427));
	DIV428: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(395), SI=>SUB_SOS(396), BI=>SUB_BOS(427), OKI=>SUB_OKOS(429), BO=>SUB_BOS(428), OKO=>SUB_OKOS(428), D=>SUB_DS(428), SO=>SUB_SOS(428));
	DIV429: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(396), SI=>SUB_SOS(397), BI=>SUB_BOS(428), OKI=>SUB_OKOS(430), BO=>SUB_BOS(429), OKO=>SUB_OKOS(429), D=>SUB_DS(429), SO=>SUB_SOS(429));
	DIV430: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(397), SI=>SUB_SOS(398), BI=>SUB_BOS(429), OKI=>SUB_OKOS(431), BO=>SUB_BOS(430), OKO=>SUB_OKOS(430), D=>SUB_DS(430), SO=>SUB_SOS(430));
	DIV431: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(398), SI=>SUB_SOS(399), BI=>SUB_BOS(430), OKI=>SUB_OKOS(432), BO=>SUB_BOS(431), OKO=>SUB_OKOS(431), D=>SUB_DS(431), SO=>SUB_SOS(431));
	DIV432: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(399), SI=>SUB_SOS(400), BI=>SUB_BOS(431), OKI=>SUB_OKOS(433), BO=>SUB_BOS(432), OKO=>SUB_OKOS(432), D=>SUB_DS(432), SO=>SUB_SOS(432));
	DIV433: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(400), SI=>SUB_SOS(401), BI=>SUB_BOS(432), OKI=>SUB_OKOS(434), BO=>SUB_BOS(433), OKO=>SUB_OKOS(433), D=>SUB_DS(433), SO=>SUB_SOS(433));
	DIV434: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(401), SI=>SUB_SOS(402), BI=>SUB_BOS(433), OKI=>SUB_OKOS(435), BO=>SUB_BOS(434), OKO=>SUB_OKOS(434), D=>SUB_DS(434), SO=>SUB_SOS(434));
	DIV435: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(402), SI=>SUB_SOS(403), BI=>SUB_BOS(434), OKI=>SUB_OKOS(436), BO=>SUB_BOS(435), OKO=>SUB_OKOS(435), D=>SUB_DS(435), SO=>SUB_SOS(435));
	DIV436: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(403), SI=>SUB_SOS(404), BI=>SUB_BOS(435), OKI=>SUB_OKOS(437), BO=>SUB_BOS(436), OKO=>SUB_OKOS(436), D=>SUB_DS(436), SO=>SUB_SOS(436));
	DIV437: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(404), SI=>SUB_SOS(405), BI=>SUB_BOS(436), OKI=>SUB_OKOS(438), BO=>SUB_BOS(437), OKO=>SUB_OKOS(437), D=>SUB_DS(437), SO=>SUB_SOS(437));
	DIV438: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(405), SI=>SUB_SOS(406), BI=>SUB_BOS(437), OKI=>SUB_OKOS(439), BO=>SUB_BOS(438), OKO=>SUB_OKOS(438), D=>SUB_DS(438), SO=>SUB_SOS(438));
	DIV439: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(406), SI=>SUB_SOS(407), BI=>SUB_BOS(438), OKI=>SUB_OKOS(440), BO=>SUB_BOS(439), OKO=>SUB_OKOS(439), D=>SUB_DS(439), SO=>SUB_SOS(439));
	DIV440: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(407), SI=>SUB_SOS(408), BI=>SUB_BOS(439), OKI=>SUB_OKOS(441), BO=>SUB_BOS(440), OKO=>SUB_OKOS(440), D=>SUB_DS(440), SO=>SUB_SOS(440));
	DIV441: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(408), SI=>SUB_SOS(409), BI=>SUB_BOS(440), OKI=>SUB_OKOS(442), BO=>SUB_BOS(441), OKO=>SUB_OKOS(441), D=>SUB_DS(441), SO=>SUB_SOS(441));
	DIV442: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(409), SI=>SUB_SOS(410), BI=>SUB_BOS(441), OKI=>SUB_OKOS(443), BO=>SUB_BOS(442), OKO=>SUB_OKOS(442), D=>SUB_DS(442), SO=>SUB_SOS(442));
	DIV443: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(410), SI=>SUB_SOS(411), BI=>SUB_BOS(442), OKI=>SUB_OKOS(444), BO=>SUB_BOS(443), OKO=>SUB_OKOS(443), D=>SUB_DS(443), SO=>SUB_SOS(443));
	DIV444: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(411), SI=>SUB_SOS(412), BI=>SUB_BOS(443), OKI=>SUB_OKOS(445), BO=>SUB_BOS(444), OKO=>SUB_OKOS(444), D=>SUB_DS(444), SO=>SUB_SOS(444));
	DIV445: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(412), SI=>SUB_SOS(413), BI=>SUB_BOS(444), OKI=>SUB_OKOS(446), BO=>SUB_BOS(445), OKO=>SUB_OKOS(445), D=>SUB_DS(445), SO=>SUB_SOS(445));
	DIV446: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(413), SI=>SUB_SOS(414), BI=>SUB_BOS(445), OKI=>SUB_OKOS(447), BO=>SUB_BOS(446), OKO=>SUB_OKOS(446), D=>SUB_DS(446), SO=>SUB_SOS(446));
	DIV447: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(414), SI=>SUB_SOS(415), BI=>SUB_BOS(446), OKI=>BONS(13), BO=>SUB_BOS(447), OKO=>SUB_OKOS(447), D=>SUB_DS(447), SO=>SUB_SOS(447));

	DIV448: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(17), SI=>SUB_SOS(416), BI=>'0', OKI=>SUB_OKOS(449), BO=>SUB_BOS(448), OKO=>SUB_OKOS(448), D=>SUB_DS(448), SO=>SUB_SOS(448));
	DIV449: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(416), SI=>SUB_SOS(417), BI=>SUB_BOS(448), OKI=>SUB_OKOS(450), BO=>SUB_BOS(449), OKO=>SUB_OKOS(449), D=>SUB_DS(449), SO=>SUB_SOS(449));
	DIV450: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(417), SI=>SUB_SOS(418), BI=>SUB_BOS(449), OKI=>SUB_OKOS(451), BO=>SUB_BOS(450), OKO=>SUB_OKOS(450), D=>SUB_DS(450), SO=>SUB_SOS(450));
	DIV451: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(418), SI=>SUB_SOS(419), BI=>SUB_BOS(450), OKI=>SUB_OKOS(452), BO=>SUB_BOS(451), OKO=>SUB_OKOS(451), D=>SUB_DS(451), SO=>SUB_SOS(451));
	DIV452: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(419), SI=>SUB_SOS(420), BI=>SUB_BOS(451), OKI=>SUB_OKOS(453), BO=>SUB_BOS(452), OKO=>SUB_OKOS(452), D=>SUB_DS(452), SO=>SUB_SOS(452));
	DIV453: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(420), SI=>SUB_SOS(421), BI=>SUB_BOS(452), OKI=>SUB_OKOS(454), BO=>SUB_BOS(453), OKO=>SUB_OKOS(453), D=>SUB_DS(453), SO=>SUB_SOS(453));
	DIV454: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(421), SI=>SUB_SOS(422), BI=>SUB_BOS(453), OKI=>SUB_OKOS(455), BO=>SUB_BOS(454), OKO=>SUB_OKOS(454), D=>SUB_DS(454), SO=>SUB_SOS(454));
	DIV455: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(422), SI=>SUB_SOS(423), BI=>SUB_BOS(454), OKI=>SUB_OKOS(456), BO=>SUB_BOS(455), OKO=>SUB_OKOS(455), D=>SUB_DS(455), SO=>SUB_SOS(455));
	DIV456: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(423), SI=>SUB_SOS(424), BI=>SUB_BOS(455), OKI=>SUB_OKOS(457), BO=>SUB_BOS(456), OKO=>SUB_OKOS(456), D=>SUB_DS(456), SO=>SUB_SOS(456));
	DIV457: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(424), SI=>SUB_SOS(425), BI=>SUB_BOS(456), OKI=>SUB_OKOS(458), BO=>SUB_BOS(457), OKO=>SUB_OKOS(457), D=>SUB_DS(457), SO=>SUB_SOS(457));
	DIV458: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(425), SI=>SUB_SOS(426), BI=>SUB_BOS(457), OKI=>SUB_OKOS(459), BO=>SUB_BOS(458), OKO=>SUB_OKOS(458), D=>SUB_DS(458), SO=>SUB_SOS(458));
	DIV459: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(426), SI=>SUB_SOS(427), BI=>SUB_BOS(458), OKI=>SUB_OKOS(460), BO=>SUB_BOS(459), OKO=>SUB_OKOS(459), D=>SUB_DS(459), SO=>SUB_SOS(459));
	DIV460: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(427), SI=>SUB_SOS(428), BI=>SUB_BOS(459), OKI=>SUB_OKOS(461), BO=>SUB_BOS(460), OKO=>SUB_OKOS(460), D=>SUB_DS(460), SO=>SUB_SOS(460));
	DIV461: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(428), SI=>SUB_SOS(429), BI=>SUB_BOS(460), OKI=>SUB_OKOS(462), BO=>SUB_BOS(461), OKO=>SUB_OKOS(461), D=>SUB_DS(461), SO=>SUB_SOS(461));
	DIV462: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(429), SI=>SUB_SOS(430), BI=>SUB_BOS(461), OKI=>SUB_OKOS(463), BO=>SUB_BOS(462), OKO=>SUB_OKOS(462), D=>SUB_DS(462), SO=>SUB_SOS(462));
	DIV463: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(430), SI=>SUB_SOS(431), BI=>SUB_BOS(462), OKI=>SUB_OKOS(464), BO=>SUB_BOS(463), OKO=>SUB_OKOS(463), D=>SUB_DS(463), SO=>SUB_SOS(463));
	DIV464: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(431), SI=>SUB_SOS(432), BI=>SUB_BOS(463), OKI=>SUB_OKOS(465), BO=>SUB_BOS(464), OKO=>SUB_OKOS(464), D=>SUB_DS(464), SO=>SUB_SOS(464));
	DIV465: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(432), SI=>SUB_SOS(433), BI=>SUB_BOS(464), OKI=>SUB_OKOS(466), BO=>SUB_BOS(465), OKO=>SUB_OKOS(465), D=>SUB_DS(465), SO=>SUB_SOS(465));
	DIV466: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(433), SI=>SUB_SOS(434), BI=>SUB_BOS(465), OKI=>SUB_OKOS(467), BO=>SUB_BOS(466), OKO=>SUB_OKOS(466), D=>SUB_DS(466), SO=>SUB_SOS(466));
	DIV467: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(434), SI=>SUB_SOS(435), BI=>SUB_BOS(466), OKI=>SUB_OKOS(468), BO=>SUB_BOS(467), OKO=>SUB_OKOS(467), D=>SUB_DS(467), SO=>SUB_SOS(467));
	DIV468: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(435), SI=>SUB_SOS(436), BI=>SUB_BOS(467), OKI=>SUB_OKOS(469), BO=>SUB_BOS(468), OKO=>SUB_OKOS(468), D=>SUB_DS(468), SO=>SUB_SOS(468));
	DIV469: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(436), SI=>SUB_SOS(437), BI=>SUB_BOS(468), OKI=>SUB_OKOS(470), BO=>SUB_BOS(469), OKO=>SUB_OKOS(469), D=>SUB_DS(469), SO=>SUB_SOS(469));
	DIV470: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(437), SI=>SUB_SOS(438), BI=>SUB_BOS(469), OKI=>SUB_OKOS(471), BO=>SUB_BOS(470), OKO=>SUB_OKOS(470), D=>SUB_DS(470), SO=>SUB_SOS(470));
	DIV471: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(438), SI=>SUB_SOS(439), BI=>SUB_BOS(470), OKI=>SUB_OKOS(472), BO=>SUB_BOS(471), OKO=>SUB_OKOS(471), D=>SUB_DS(471), SO=>SUB_SOS(471));
	DIV472: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(439), SI=>SUB_SOS(440), BI=>SUB_BOS(471), OKI=>SUB_OKOS(473), BO=>SUB_BOS(472), OKO=>SUB_OKOS(472), D=>SUB_DS(472), SO=>SUB_SOS(472));
	DIV473: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(440), SI=>SUB_SOS(441), BI=>SUB_BOS(472), OKI=>SUB_OKOS(474), BO=>SUB_BOS(473), OKO=>SUB_OKOS(473), D=>SUB_DS(473), SO=>SUB_SOS(473));
	DIV474: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(441), SI=>SUB_SOS(442), BI=>SUB_BOS(473), OKI=>SUB_OKOS(475), BO=>SUB_BOS(474), OKO=>SUB_OKOS(474), D=>SUB_DS(474), SO=>SUB_SOS(474));
	DIV475: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(442), SI=>SUB_SOS(443), BI=>SUB_BOS(474), OKI=>SUB_OKOS(476), BO=>SUB_BOS(475), OKO=>SUB_OKOS(475), D=>SUB_DS(475), SO=>SUB_SOS(475));
	DIV476: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(443), SI=>SUB_SOS(444), BI=>SUB_BOS(475), OKI=>SUB_OKOS(477), BO=>SUB_BOS(476), OKO=>SUB_OKOS(476), D=>SUB_DS(476), SO=>SUB_SOS(476));
	DIV477: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(444), SI=>SUB_SOS(445), BI=>SUB_BOS(476), OKI=>SUB_OKOS(478), BO=>SUB_BOS(477), OKO=>SUB_OKOS(477), D=>SUB_DS(477), SO=>SUB_SOS(477));
	DIV478: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(445), SI=>SUB_SOS(446), BI=>SUB_BOS(477), OKI=>SUB_OKOS(479), BO=>SUB_BOS(478), OKO=>SUB_OKOS(478), D=>SUB_DS(478), SO=>SUB_SOS(478));
	DIV479: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(446), SI=>SUB_SOS(447), BI=>SUB_BOS(478), OKI=>BONS(14), BO=>SUB_BOS(479), OKO=>SUB_OKOS(479), D=>SUB_DS(479), SO=>SUB_SOS(479));

	DIV480: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(16), SI=>SUB_SOS(448), BI=>'0', OKI=>SUB_OKOS(481), BO=>SUB_BOS(480), OKO=>SUB_OKOS(480), D=>SUB_DS(480), SO=>SUB_SOS(480));
	DIV481: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(448), SI=>SUB_SOS(449), BI=>SUB_BOS(480), OKI=>SUB_OKOS(482), BO=>SUB_BOS(481), OKO=>SUB_OKOS(481), D=>SUB_DS(481), SO=>SUB_SOS(481));
	DIV482: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(449), SI=>SUB_SOS(450), BI=>SUB_BOS(481), OKI=>SUB_OKOS(483), BO=>SUB_BOS(482), OKO=>SUB_OKOS(482), D=>SUB_DS(482), SO=>SUB_SOS(482));
	DIV483: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(450), SI=>SUB_SOS(451), BI=>SUB_BOS(482), OKI=>SUB_OKOS(484), BO=>SUB_BOS(483), OKO=>SUB_OKOS(483), D=>SUB_DS(483), SO=>SUB_SOS(483));
	DIV484: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(451), SI=>SUB_SOS(452), BI=>SUB_BOS(483), OKI=>SUB_OKOS(485), BO=>SUB_BOS(484), OKO=>SUB_OKOS(484), D=>SUB_DS(484), SO=>SUB_SOS(484));
	DIV485: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(452), SI=>SUB_SOS(453), BI=>SUB_BOS(484), OKI=>SUB_OKOS(486), BO=>SUB_BOS(485), OKO=>SUB_OKOS(485), D=>SUB_DS(485), SO=>SUB_SOS(485));
	DIV486: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(453), SI=>SUB_SOS(454), BI=>SUB_BOS(485), OKI=>SUB_OKOS(487), BO=>SUB_BOS(486), OKO=>SUB_OKOS(486), D=>SUB_DS(486), SO=>SUB_SOS(486));
	DIV487: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(454), SI=>SUB_SOS(455), BI=>SUB_BOS(486), OKI=>SUB_OKOS(488), BO=>SUB_BOS(487), OKO=>SUB_OKOS(487), D=>SUB_DS(487), SO=>SUB_SOS(487));
	DIV488: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(455), SI=>SUB_SOS(456), BI=>SUB_BOS(487), OKI=>SUB_OKOS(489), BO=>SUB_BOS(488), OKO=>SUB_OKOS(488), D=>SUB_DS(488), SO=>SUB_SOS(488));
	DIV489: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(456), SI=>SUB_SOS(457), BI=>SUB_BOS(488), OKI=>SUB_OKOS(490), BO=>SUB_BOS(489), OKO=>SUB_OKOS(489), D=>SUB_DS(489), SO=>SUB_SOS(489));
	DIV490: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(457), SI=>SUB_SOS(458), BI=>SUB_BOS(489), OKI=>SUB_OKOS(491), BO=>SUB_BOS(490), OKO=>SUB_OKOS(490), D=>SUB_DS(490), SO=>SUB_SOS(490));
	DIV491: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(458), SI=>SUB_SOS(459), BI=>SUB_BOS(490), OKI=>SUB_OKOS(492), BO=>SUB_BOS(491), OKO=>SUB_OKOS(491), D=>SUB_DS(491), SO=>SUB_SOS(491));
	DIV492: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(459), SI=>SUB_SOS(460), BI=>SUB_BOS(491), OKI=>SUB_OKOS(493), BO=>SUB_BOS(492), OKO=>SUB_OKOS(492), D=>SUB_DS(492), SO=>SUB_SOS(492));
	DIV493: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(460), SI=>SUB_SOS(461), BI=>SUB_BOS(492), OKI=>SUB_OKOS(494), BO=>SUB_BOS(493), OKO=>SUB_OKOS(493), D=>SUB_DS(493), SO=>SUB_SOS(493));
	DIV494: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(461), SI=>SUB_SOS(462), BI=>SUB_BOS(493), OKI=>SUB_OKOS(495), BO=>SUB_BOS(494), OKO=>SUB_OKOS(494), D=>SUB_DS(494), SO=>SUB_SOS(494));
	DIV495: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(462), SI=>SUB_SOS(463), BI=>SUB_BOS(494), OKI=>SUB_OKOS(496), BO=>SUB_BOS(495), OKO=>SUB_OKOS(495), D=>SUB_DS(495), SO=>SUB_SOS(495));
	DIV496: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(463), SI=>SUB_SOS(464), BI=>SUB_BOS(495), OKI=>SUB_OKOS(497), BO=>SUB_BOS(496), OKO=>SUB_OKOS(496), D=>SUB_DS(496), SO=>SUB_SOS(496));
	DIV497: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(464), SI=>SUB_SOS(465), BI=>SUB_BOS(496), OKI=>SUB_OKOS(498), BO=>SUB_BOS(497), OKO=>SUB_OKOS(497), D=>SUB_DS(497), SO=>SUB_SOS(497));
	DIV498: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(465), SI=>SUB_SOS(466), BI=>SUB_BOS(497), OKI=>SUB_OKOS(499), BO=>SUB_BOS(498), OKO=>SUB_OKOS(498), D=>SUB_DS(498), SO=>SUB_SOS(498));
	DIV499: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(466), SI=>SUB_SOS(467), BI=>SUB_BOS(498), OKI=>SUB_OKOS(500), BO=>SUB_BOS(499), OKO=>SUB_OKOS(499), D=>SUB_DS(499), SO=>SUB_SOS(499));
	DIV500: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(467), SI=>SUB_SOS(468), BI=>SUB_BOS(499), OKI=>SUB_OKOS(501), BO=>SUB_BOS(500), OKO=>SUB_OKOS(500), D=>SUB_DS(500), SO=>SUB_SOS(500));
	DIV501: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(468), SI=>SUB_SOS(469), BI=>SUB_BOS(500), OKI=>SUB_OKOS(502), BO=>SUB_BOS(501), OKO=>SUB_OKOS(501), D=>SUB_DS(501), SO=>SUB_SOS(501));
	DIV502: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(469), SI=>SUB_SOS(470), BI=>SUB_BOS(501), OKI=>SUB_OKOS(503), BO=>SUB_BOS(502), OKO=>SUB_OKOS(502), D=>SUB_DS(502), SO=>SUB_SOS(502));
	DIV503: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(470), SI=>SUB_SOS(471), BI=>SUB_BOS(502), OKI=>SUB_OKOS(504), BO=>SUB_BOS(503), OKO=>SUB_OKOS(503), D=>SUB_DS(503), SO=>SUB_SOS(503));
	DIV504: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(471), SI=>SUB_SOS(472), BI=>SUB_BOS(503), OKI=>SUB_OKOS(505), BO=>SUB_BOS(504), OKO=>SUB_OKOS(504), D=>SUB_DS(504), SO=>SUB_SOS(504));
	DIV505: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(472), SI=>SUB_SOS(473), BI=>SUB_BOS(504), OKI=>SUB_OKOS(506), BO=>SUB_BOS(505), OKO=>SUB_OKOS(505), D=>SUB_DS(505), SO=>SUB_SOS(505));
	DIV506: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(473), SI=>SUB_SOS(474), BI=>SUB_BOS(505), OKI=>SUB_OKOS(507), BO=>SUB_BOS(506), OKO=>SUB_OKOS(506), D=>SUB_DS(506), SO=>SUB_SOS(506));
	DIV507: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(474), SI=>SUB_SOS(475), BI=>SUB_BOS(506), OKI=>SUB_OKOS(508), BO=>SUB_BOS(507), OKO=>SUB_OKOS(507), D=>SUB_DS(507), SO=>SUB_SOS(507));
	DIV508: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(475), SI=>SUB_SOS(476), BI=>SUB_BOS(507), OKI=>SUB_OKOS(509), BO=>SUB_BOS(508), OKO=>SUB_OKOS(508), D=>SUB_DS(508), SO=>SUB_SOS(508));
	DIV509: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(476), SI=>SUB_SOS(477), BI=>SUB_BOS(508), OKI=>SUB_OKOS(510), BO=>SUB_BOS(509), OKO=>SUB_OKOS(509), D=>SUB_DS(509), SO=>SUB_SOS(509));
	DIV510: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(477), SI=>SUB_SOS(478), BI=>SUB_BOS(509), OKI=>SUB_OKOS(511), BO=>SUB_BOS(510), OKO=>SUB_OKOS(510), D=>SUB_DS(510), SO=>SUB_SOS(510));
	DIV511: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(478), SI=>SUB_SOS(479), BI=>SUB_BOS(510), OKI=>BONS(15), BO=>SUB_BOS(511), OKO=>SUB_OKOS(511), D=>SUB_DS(511), SO=>SUB_SOS(511));

	DIV512: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(15), SI=>SUB_SOS(480), BI=>'0', OKI=>SUB_OKOS(513), BO=>SUB_BOS(512), OKO=>SUB_OKOS(512), D=>SUB_DS(512), SO=>SUB_SOS(512));
	DIV513: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(480), SI=>SUB_SOS(481), BI=>SUB_BOS(512), OKI=>SUB_OKOS(514), BO=>SUB_BOS(513), OKO=>SUB_OKOS(513), D=>SUB_DS(513), SO=>SUB_SOS(513));
	DIV514: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(481), SI=>SUB_SOS(482), BI=>SUB_BOS(513), OKI=>SUB_OKOS(515), BO=>SUB_BOS(514), OKO=>SUB_OKOS(514), D=>SUB_DS(514), SO=>SUB_SOS(514));
	DIV515: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(482), SI=>SUB_SOS(483), BI=>SUB_BOS(514), OKI=>SUB_OKOS(516), BO=>SUB_BOS(515), OKO=>SUB_OKOS(515), D=>SUB_DS(515), SO=>SUB_SOS(515));
	DIV516: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(483), SI=>SUB_SOS(484), BI=>SUB_BOS(515), OKI=>SUB_OKOS(517), BO=>SUB_BOS(516), OKO=>SUB_OKOS(516), D=>SUB_DS(516), SO=>SUB_SOS(516));
	DIV517: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(484), SI=>SUB_SOS(485), BI=>SUB_BOS(516), OKI=>SUB_OKOS(518), BO=>SUB_BOS(517), OKO=>SUB_OKOS(517), D=>SUB_DS(517), SO=>SUB_SOS(517));
	DIV518: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(485), SI=>SUB_SOS(486), BI=>SUB_BOS(517), OKI=>SUB_OKOS(519), BO=>SUB_BOS(518), OKO=>SUB_OKOS(518), D=>SUB_DS(518), SO=>SUB_SOS(518));
	DIV519: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(486), SI=>SUB_SOS(487), BI=>SUB_BOS(518), OKI=>SUB_OKOS(520), BO=>SUB_BOS(519), OKO=>SUB_OKOS(519), D=>SUB_DS(519), SO=>SUB_SOS(519));
	DIV520: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(487), SI=>SUB_SOS(488), BI=>SUB_BOS(519), OKI=>SUB_OKOS(521), BO=>SUB_BOS(520), OKO=>SUB_OKOS(520), D=>SUB_DS(520), SO=>SUB_SOS(520));
	DIV521: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(488), SI=>SUB_SOS(489), BI=>SUB_BOS(520), OKI=>SUB_OKOS(522), BO=>SUB_BOS(521), OKO=>SUB_OKOS(521), D=>SUB_DS(521), SO=>SUB_SOS(521));
	DIV522: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(489), SI=>SUB_SOS(490), BI=>SUB_BOS(521), OKI=>SUB_OKOS(523), BO=>SUB_BOS(522), OKO=>SUB_OKOS(522), D=>SUB_DS(522), SO=>SUB_SOS(522));
	DIV523: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(490), SI=>SUB_SOS(491), BI=>SUB_BOS(522), OKI=>SUB_OKOS(524), BO=>SUB_BOS(523), OKO=>SUB_OKOS(523), D=>SUB_DS(523), SO=>SUB_SOS(523));
	DIV524: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(491), SI=>SUB_SOS(492), BI=>SUB_BOS(523), OKI=>SUB_OKOS(525), BO=>SUB_BOS(524), OKO=>SUB_OKOS(524), D=>SUB_DS(524), SO=>SUB_SOS(524));
	DIV525: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(492), SI=>SUB_SOS(493), BI=>SUB_BOS(524), OKI=>SUB_OKOS(526), BO=>SUB_BOS(525), OKO=>SUB_OKOS(525), D=>SUB_DS(525), SO=>SUB_SOS(525));
	DIV526: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(493), SI=>SUB_SOS(494), BI=>SUB_BOS(525), OKI=>SUB_OKOS(527), BO=>SUB_BOS(526), OKO=>SUB_OKOS(526), D=>SUB_DS(526), SO=>SUB_SOS(526));
	DIV527: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(494), SI=>SUB_SOS(495), BI=>SUB_BOS(526), OKI=>SUB_OKOS(528), BO=>SUB_BOS(527), OKO=>SUB_OKOS(527), D=>SUB_DS(527), SO=>SUB_SOS(527));
	DIV528: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(495), SI=>SUB_SOS(496), BI=>SUB_BOS(527), OKI=>SUB_OKOS(529), BO=>SUB_BOS(528), OKO=>SUB_OKOS(528), D=>SUB_DS(528), SO=>SUB_SOS(528));
	DIV529: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(496), SI=>SUB_SOS(497), BI=>SUB_BOS(528), OKI=>SUB_OKOS(530), BO=>SUB_BOS(529), OKO=>SUB_OKOS(529), D=>SUB_DS(529), SO=>SUB_SOS(529));
	DIV530: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(497), SI=>SUB_SOS(498), BI=>SUB_BOS(529), OKI=>SUB_OKOS(531), BO=>SUB_BOS(530), OKO=>SUB_OKOS(530), D=>SUB_DS(530), SO=>SUB_SOS(530));
	DIV531: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(498), SI=>SUB_SOS(499), BI=>SUB_BOS(530), OKI=>SUB_OKOS(532), BO=>SUB_BOS(531), OKO=>SUB_OKOS(531), D=>SUB_DS(531), SO=>SUB_SOS(531));
	DIV532: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(499), SI=>SUB_SOS(500), BI=>SUB_BOS(531), OKI=>SUB_OKOS(533), BO=>SUB_BOS(532), OKO=>SUB_OKOS(532), D=>SUB_DS(532), SO=>SUB_SOS(532));
	DIV533: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(500), SI=>SUB_SOS(501), BI=>SUB_BOS(532), OKI=>SUB_OKOS(534), BO=>SUB_BOS(533), OKO=>SUB_OKOS(533), D=>SUB_DS(533), SO=>SUB_SOS(533));
	DIV534: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(501), SI=>SUB_SOS(502), BI=>SUB_BOS(533), OKI=>SUB_OKOS(535), BO=>SUB_BOS(534), OKO=>SUB_OKOS(534), D=>SUB_DS(534), SO=>SUB_SOS(534));
	DIV535: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(502), SI=>SUB_SOS(503), BI=>SUB_BOS(534), OKI=>SUB_OKOS(536), BO=>SUB_BOS(535), OKO=>SUB_OKOS(535), D=>SUB_DS(535), SO=>SUB_SOS(535));
	DIV536: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(503), SI=>SUB_SOS(504), BI=>SUB_BOS(535), OKI=>SUB_OKOS(537), BO=>SUB_BOS(536), OKO=>SUB_OKOS(536), D=>SUB_DS(536), SO=>SUB_SOS(536));
	DIV537: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(504), SI=>SUB_SOS(505), BI=>SUB_BOS(536), OKI=>SUB_OKOS(538), BO=>SUB_BOS(537), OKO=>SUB_OKOS(537), D=>SUB_DS(537), SO=>SUB_SOS(537));
	DIV538: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(505), SI=>SUB_SOS(506), BI=>SUB_BOS(537), OKI=>SUB_OKOS(539), BO=>SUB_BOS(538), OKO=>SUB_OKOS(538), D=>SUB_DS(538), SO=>SUB_SOS(538));
	DIV539: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(506), SI=>SUB_SOS(507), BI=>SUB_BOS(538), OKI=>SUB_OKOS(540), BO=>SUB_BOS(539), OKO=>SUB_OKOS(539), D=>SUB_DS(539), SO=>SUB_SOS(539));
	DIV540: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(507), SI=>SUB_SOS(508), BI=>SUB_BOS(539), OKI=>SUB_OKOS(541), BO=>SUB_BOS(540), OKO=>SUB_OKOS(540), D=>SUB_DS(540), SO=>SUB_SOS(540));
	DIV541: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(508), SI=>SUB_SOS(509), BI=>SUB_BOS(540), OKI=>SUB_OKOS(542), BO=>SUB_BOS(541), OKO=>SUB_OKOS(541), D=>SUB_DS(541), SO=>SUB_SOS(541));
	DIV542: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(509), SI=>SUB_SOS(510), BI=>SUB_BOS(541), OKI=>SUB_OKOS(543), BO=>SUB_BOS(542), OKO=>SUB_OKOS(542), D=>SUB_DS(542), SO=>SUB_SOS(542));
	DIV543: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(510), SI=>SUB_SOS(511), BI=>SUB_BOS(542), OKI=>BONS(16), BO=>SUB_BOS(543), OKO=>SUB_OKOS(543), D=>SUB_DS(543), SO=>SUB_SOS(543));

	DIV544: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(14), SI=>SUB_SOS(512), BI=>'0', OKI=>SUB_OKOS(545), BO=>SUB_BOS(544), OKO=>SUB_OKOS(544), D=>SUB_DS(544), SO=>SUB_SOS(544));
	DIV545: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(512), SI=>SUB_SOS(513), BI=>SUB_BOS(544), OKI=>SUB_OKOS(546), BO=>SUB_BOS(545), OKO=>SUB_OKOS(545), D=>SUB_DS(545), SO=>SUB_SOS(545));
	DIV546: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(513), SI=>SUB_SOS(514), BI=>SUB_BOS(545), OKI=>SUB_OKOS(547), BO=>SUB_BOS(546), OKO=>SUB_OKOS(546), D=>SUB_DS(546), SO=>SUB_SOS(546));
	DIV547: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(514), SI=>SUB_SOS(515), BI=>SUB_BOS(546), OKI=>SUB_OKOS(548), BO=>SUB_BOS(547), OKO=>SUB_OKOS(547), D=>SUB_DS(547), SO=>SUB_SOS(547));
	DIV548: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(515), SI=>SUB_SOS(516), BI=>SUB_BOS(547), OKI=>SUB_OKOS(549), BO=>SUB_BOS(548), OKO=>SUB_OKOS(548), D=>SUB_DS(548), SO=>SUB_SOS(548));
	DIV549: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(516), SI=>SUB_SOS(517), BI=>SUB_BOS(548), OKI=>SUB_OKOS(550), BO=>SUB_BOS(549), OKO=>SUB_OKOS(549), D=>SUB_DS(549), SO=>SUB_SOS(549));
	DIV550: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(517), SI=>SUB_SOS(518), BI=>SUB_BOS(549), OKI=>SUB_OKOS(551), BO=>SUB_BOS(550), OKO=>SUB_OKOS(550), D=>SUB_DS(550), SO=>SUB_SOS(550));
	DIV551: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(518), SI=>SUB_SOS(519), BI=>SUB_BOS(550), OKI=>SUB_OKOS(552), BO=>SUB_BOS(551), OKO=>SUB_OKOS(551), D=>SUB_DS(551), SO=>SUB_SOS(551));
	DIV552: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(519), SI=>SUB_SOS(520), BI=>SUB_BOS(551), OKI=>SUB_OKOS(553), BO=>SUB_BOS(552), OKO=>SUB_OKOS(552), D=>SUB_DS(552), SO=>SUB_SOS(552));
	DIV553: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(520), SI=>SUB_SOS(521), BI=>SUB_BOS(552), OKI=>SUB_OKOS(554), BO=>SUB_BOS(553), OKO=>SUB_OKOS(553), D=>SUB_DS(553), SO=>SUB_SOS(553));
	DIV554: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(521), SI=>SUB_SOS(522), BI=>SUB_BOS(553), OKI=>SUB_OKOS(555), BO=>SUB_BOS(554), OKO=>SUB_OKOS(554), D=>SUB_DS(554), SO=>SUB_SOS(554));
	DIV555: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(522), SI=>SUB_SOS(523), BI=>SUB_BOS(554), OKI=>SUB_OKOS(556), BO=>SUB_BOS(555), OKO=>SUB_OKOS(555), D=>SUB_DS(555), SO=>SUB_SOS(555));
	DIV556: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(523), SI=>SUB_SOS(524), BI=>SUB_BOS(555), OKI=>SUB_OKOS(557), BO=>SUB_BOS(556), OKO=>SUB_OKOS(556), D=>SUB_DS(556), SO=>SUB_SOS(556));
	DIV557: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(524), SI=>SUB_SOS(525), BI=>SUB_BOS(556), OKI=>SUB_OKOS(558), BO=>SUB_BOS(557), OKO=>SUB_OKOS(557), D=>SUB_DS(557), SO=>SUB_SOS(557));
	DIV558: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(525), SI=>SUB_SOS(526), BI=>SUB_BOS(557), OKI=>SUB_OKOS(559), BO=>SUB_BOS(558), OKO=>SUB_OKOS(558), D=>SUB_DS(558), SO=>SUB_SOS(558));
	DIV559: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(526), SI=>SUB_SOS(527), BI=>SUB_BOS(558), OKI=>SUB_OKOS(560), BO=>SUB_BOS(559), OKO=>SUB_OKOS(559), D=>SUB_DS(559), SO=>SUB_SOS(559));
	DIV560: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(527), SI=>SUB_SOS(528), BI=>SUB_BOS(559), OKI=>SUB_OKOS(561), BO=>SUB_BOS(560), OKO=>SUB_OKOS(560), D=>SUB_DS(560), SO=>SUB_SOS(560));
	DIV561: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(528), SI=>SUB_SOS(529), BI=>SUB_BOS(560), OKI=>SUB_OKOS(562), BO=>SUB_BOS(561), OKO=>SUB_OKOS(561), D=>SUB_DS(561), SO=>SUB_SOS(561));
	DIV562: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(529), SI=>SUB_SOS(530), BI=>SUB_BOS(561), OKI=>SUB_OKOS(563), BO=>SUB_BOS(562), OKO=>SUB_OKOS(562), D=>SUB_DS(562), SO=>SUB_SOS(562));
	DIV563: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(530), SI=>SUB_SOS(531), BI=>SUB_BOS(562), OKI=>SUB_OKOS(564), BO=>SUB_BOS(563), OKO=>SUB_OKOS(563), D=>SUB_DS(563), SO=>SUB_SOS(563));
	DIV564: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(531), SI=>SUB_SOS(532), BI=>SUB_BOS(563), OKI=>SUB_OKOS(565), BO=>SUB_BOS(564), OKO=>SUB_OKOS(564), D=>SUB_DS(564), SO=>SUB_SOS(564));
	DIV565: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(532), SI=>SUB_SOS(533), BI=>SUB_BOS(564), OKI=>SUB_OKOS(566), BO=>SUB_BOS(565), OKO=>SUB_OKOS(565), D=>SUB_DS(565), SO=>SUB_SOS(565));
	DIV566: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(533), SI=>SUB_SOS(534), BI=>SUB_BOS(565), OKI=>SUB_OKOS(567), BO=>SUB_BOS(566), OKO=>SUB_OKOS(566), D=>SUB_DS(566), SO=>SUB_SOS(566));
	DIV567: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(534), SI=>SUB_SOS(535), BI=>SUB_BOS(566), OKI=>SUB_OKOS(568), BO=>SUB_BOS(567), OKO=>SUB_OKOS(567), D=>SUB_DS(567), SO=>SUB_SOS(567));
	DIV568: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(535), SI=>SUB_SOS(536), BI=>SUB_BOS(567), OKI=>SUB_OKOS(569), BO=>SUB_BOS(568), OKO=>SUB_OKOS(568), D=>SUB_DS(568), SO=>SUB_SOS(568));
	DIV569: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(536), SI=>SUB_SOS(537), BI=>SUB_BOS(568), OKI=>SUB_OKOS(570), BO=>SUB_BOS(569), OKO=>SUB_OKOS(569), D=>SUB_DS(569), SO=>SUB_SOS(569));
	DIV570: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(537), SI=>SUB_SOS(538), BI=>SUB_BOS(569), OKI=>SUB_OKOS(571), BO=>SUB_BOS(570), OKO=>SUB_OKOS(570), D=>SUB_DS(570), SO=>SUB_SOS(570));
	DIV571: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(538), SI=>SUB_SOS(539), BI=>SUB_BOS(570), OKI=>SUB_OKOS(572), BO=>SUB_BOS(571), OKO=>SUB_OKOS(571), D=>SUB_DS(571), SO=>SUB_SOS(571));
	DIV572: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(539), SI=>SUB_SOS(540), BI=>SUB_BOS(571), OKI=>SUB_OKOS(573), BO=>SUB_BOS(572), OKO=>SUB_OKOS(572), D=>SUB_DS(572), SO=>SUB_SOS(572));
	DIV573: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(540), SI=>SUB_SOS(541), BI=>SUB_BOS(572), OKI=>SUB_OKOS(574), BO=>SUB_BOS(573), OKO=>SUB_OKOS(573), D=>SUB_DS(573), SO=>SUB_SOS(573));
	DIV574: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(541), SI=>SUB_SOS(542), BI=>SUB_BOS(573), OKI=>SUB_OKOS(575), BO=>SUB_BOS(574), OKO=>SUB_OKOS(574), D=>SUB_DS(574), SO=>SUB_SOS(574));
	DIV575: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(542), SI=>SUB_SOS(543), BI=>SUB_BOS(574), OKI=>BONS(17), BO=>SUB_BOS(575), OKO=>SUB_OKOS(575), D=>SUB_DS(575), SO=>SUB_SOS(575));

	DIV576: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(13), SI=>SUB_SOS(544), BI=>'0', OKI=>SUB_OKOS(577), BO=>SUB_BOS(576), OKO=>SUB_OKOS(576), D=>SUB_DS(576), SO=>SUB_SOS(576));
	DIV577: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(544), SI=>SUB_SOS(545), BI=>SUB_BOS(576), OKI=>SUB_OKOS(578), BO=>SUB_BOS(577), OKO=>SUB_OKOS(577), D=>SUB_DS(577), SO=>SUB_SOS(577));
	DIV578: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(545), SI=>SUB_SOS(546), BI=>SUB_BOS(577), OKI=>SUB_OKOS(579), BO=>SUB_BOS(578), OKO=>SUB_OKOS(578), D=>SUB_DS(578), SO=>SUB_SOS(578));
	DIV579: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(546), SI=>SUB_SOS(547), BI=>SUB_BOS(578), OKI=>SUB_OKOS(580), BO=>SUB_BOS(579), OKO=>SUB_OKOS(579), D=>SUB_DS(579), SO=>SUB_SOS(579));
	DIV580: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(547), SI=>SUB_SOS(548), BI=>SUB_BOS(579), OKI=>SUB_OKOS(581), BO=>SUB_BOS(580), OKO=>SUB_OKOS(580), D=>SUB_DS(580), SO=>SUB_SOS(580));
	DIV581: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(548), SI=>SUB_SOS(549), BI=>SUB_BOS(580), OKI=>SUB_OKOS(582), BO=>SUB_BOS(581), OKO=>SUB_OKOS(581), D=>SUB_DS(581), SO=>SUB_SOS(581));
	DIV582: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(549), SI=>SUB_SOS(550), BI=>SUB_BOS(581), OKI=>SUB_OKOS(583), BO=>SUB_BOS(582), OKO=>SUB_OKOS(582), D=>SUB_DS(582), SO=>SUB_SOS(582));
	DIV583: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(550), SI=>SUB_SOS(551), BI=>SUB_BOS(582), OKI=>SUB_OKOS(584), BO=>SUB_BOS(583), OKO=>SUB_OKOS(583), D=>SUB_DS(583), SO=>SUB_SOS(583));
	DIV584: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(551), SI=>SUB_SOS(552), BI=>SUB_BOS(583), OKI=>SUB_OKOS(585), BO=>SUB_BOS(584), OKO=>SUB_OKOS(584), D=>SUB_DS(584), SO=>SUB_SOS(584));
	DIV585: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(552), SI=>SUB_SOS(553), BI=>SUB_BOS(584), OKI=>SUB_OKOS(586), BO=>SUB_BOS(585), OKO=>SUB_OKOS(585), D=>SUB_DS(585), SO=>SUB_SOS(585));
	DIV586: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(553), SI=>SUB_SOS(554), BI=>SUB_BOS(585), OKI=>SUB_OKOS(587), BO=>SUB_BOS(586), OKO=>SUB_OKOS(586), D=>SUB_DS(586), SO=>SUB_SOS(586));
	DIV587: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(554), SI=>SUB_SOS(555), BI=>SUB_BOS(586), OKI=>SUB_OKOS(588), BO=>SUB_BOS(587), OKO=>SUB_OKOS(587), D=>SUB_DS(587), SO=>SUB_SOS(587));
	DIV588: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(555), SI=>SUB_SOS(556), BI=>SUB_BOS(587), OKI=>SUB_OKOS(589), BO=>SUB_BOS(588), OKO=>SUB_OKOS(588), D=>SUB_DS(588), SO=>SUB_SOS(588));
	DIV589: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(556), SI=>SUB_SOS(557), BI=>SUB_BOS(588), OKI=>SUB_OKOS(590), BO=>SUB_BOS(589), OKO=>SUB_OKOS(589), D=>SUB_DS(589), SO=>SUB_SOS(589));
	DIV590: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(557), SI=>SUB_SOS(558), BI=>SUB_BOS(589), OKI=>SUB_OKOS(591), BO=>SUB_BOS(590), OKO=>SUB_OKOS(590), D=>SUB_DS(590), SO=>SUB_SOS(590));
	DIV591: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(558), SI=>SUB_SOS(559), BI=>SUB_BOS(590), OKI=>SUB_OKOS(592), BO=>SUB_BOS(591), OKO=>SUB_OKOS(591), D=>SUB_DS(591), SO=>SUB_SOS(591));
	DIV592: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(559), SI=>SUB_SOS(560), BI=>SUB_BOS(591), OKI=>SUB_OKOS(593), BO=>SUB_BOS(592), OKO=>SUB_OKOS(592), D=>SUB_DS(592), SO=>SUB_SOS(592));
	DIV593: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(560), SI=>SUB_SOS(561), BI=>SUB_BOS(592), OKI=>SUB_OKOS(594), BO=>SUB_BOS(593), OKO=>SUB_OKOS(593), D=>SUB_DS(593), SO=>SUB_SOS(593));
	DIV594: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(561), SI=>SUB_SOS(562), BI=>SUB_BOS(593), OKI=>SUB_OKOS(595), BO=>SUB_BOS(594), OKO=>SUB_OKOS(594), D=>SUB_DS(594), SO=>SUB_SOS(594));
	DIV595: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(562), SI=>SUB_SOS(563), BI=>SUB_BOS(594), OKI=>SUB_OKOS(596), BO=>SUB_BOS(595), OKO=>SUB_OKOS(595), D=>SUB_DS(595), SO=>SUB_SOS(595));
	DIV596: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(563), SI=>SUB_SOS(564), BI=>SUB_BOS(595), OKI=>SUB_OKOS(597), BO=>SUB_BOS(596), OKO=>SUB_OKOS(596), D=>SUB_DS(596), SO=>SUB_SOS(596));
	DIV597: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(564), SI=>SUB_SOS(565), BI=>SUB_BOS(596), OKI=>SUB_OKOS(598), BO=>SUB_BOS(597), OKO=>SUB_OKOS(597), D=>SUB_DS(597), SO=>SUB_SOS(597));
	DIV598: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(565), SI=>SUB_SOS(566), BI=>SUB_BOS(597), OKI=>SUB_OKOS(599), BO=>SUB_BOS(598), OKO=>SUB_OKOS(598), D=>SUB_DS(598), SO=>SUB_SOS(598));
	DIV599: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(566), SI=>SUB_SOS(567), BI=>SUB_BOS(598), OKI=>SUB_OKOS(600), BO=>SUB_BOS(599), OKO=>SUB_OKOS(599), D=>SUB_DS(599), SO=>SUB_SOS(599));
	DIV600: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(567), SI=>SUB_SOS(568), BI=>SUB_BOS(599), OKI=>SUB_OKOS(601), BO=>SUB_BOS(600), OKO=>SUB_OKOS(600), D=>SUB_DS(600), SO=>SUB_SOS(600));
	DIV601: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(568), SI=>SUB_SOS(569), BI=>SUB_BOS(600), OKI=>SUB_OKOS(602), BO=>SUB_BOS(601), OKO=>SUB_OKOS(601), D=>SUB_DS(601), SO=>SUB_SOS(601));
	DIV602: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(569), SI=>SUB_SOS(570), BI=>SUB_BOS(601), OKI=>SUB_OKOS(603), BO=>SUB_BOS(602), OKO=>SUB_OKOS(602), D=>SUB_DS(602), SO=>SUB_SOS(602));
	DIV603: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(570), SI=>SUB_SOS(571), BI=>SUB_BOS(602), OKI=>SUB_OKOS(604), BO=>SUB_BOS(603), OKO=>SUB_OKOS(603), D=>SUB_DS(603), SO=>SUB_SOS(603));
	DIV604: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(571), SI=>SUB_SOS(572), BI=>SUB_BOS(603), OKI=>SUB_OKOS(605), BO=>SUB_BOS(604), OKO=>SUB_OKOS(604), D=>SUB_DS(604), SO=>SUB_SOS(604));
	DIV605: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(572), SI=>SUB_SOS(573), BI=>SUB_BOS(604), OKI=>SUB_OKOS(606), BO=>SUB_BOS(605), OKO=>SUB_OKOS(605), D=>SUB_DS(605), SO=>SUB_SOS(605));
	DIV606: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(573), SI=>SUB_SOS(574), BI=>SUB_BOS(605), OKI=>SUB_OKOS(607), BO=>SUB_BOS(606), OKO=>SUB_OKOS(606), D=>SUB_DS(606), SO=>SUB_SOS(606));
	DIV607: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(574), SI=>SUB_SOS(575), BI=>SUB_BOS(606), OKI=>BONS(18), BO=>SUB_BOS(607), OKO=>SUB_OKOS(607), D=>SUB_DS(607), SO=>SUB_SOS(607));

	DIV608: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(12), SI=>SUB_SOS(576), BI=>'0', OKI=>SUB_OKOS(609), BO=>SUB_BOS(608), OKO=>SUB_OKOS(608), D=>SUB_DS(608), SO=>SUB_SOS(608));
	DIV609: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(576), SI=>SUB_SOS(577), BI=>SUB_BOS(608), OKI=>SUB_OKOS(610), BO=>SUB_BOS(609), OKO=>SUB_OKOS(609), D=>SUB_DS(609), SO=>SUB_SOS(609));
	DIV610: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(577), SI=>SUB_SOS(578), BI=>SUB_BOS(609), OKI=>SUB_OKOS(611), BO=>SUB_BOS(610), OKO=>SUB_OKOS(610), D=>SUB_DS(610), SO=>SUB_SOS(610));
	DIV611: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(578), SI=>SUB_SOS(579), BI=>SUB_BOS(610), OKI=>SUB_OKOS(612), BO=>SUB_BOS(611), OKO=>SUB_OKOS(611), D=>SUB_DS(611), SO=>SUB_SOS(611));
	DIV612: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(579), SI=>SUB_SOS(580), BI=>SUB_BOS(611), OKI=>SUB_OKOS(613), BO=>SUB_BOS(612), OKO=>SUB_OKOS(612), D=>SUB_DS(612), SO=>SUB_SOS(612));
	DIV613: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(580), SI=>SUB_SOS(581), BI=>SUB_BOS(612), OKI=>SUB_OKOS(614), BO=>SUB_BOS(613), OKO=>SUB_OKOS(613), D=>SUB_DS(613), SO=>SUB_SOS(613));
	DIV614: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(581), SI=>SUB_SOS(582), BI=>SUB_BOS(613), OKI=>SUB_OKOS(615), BO=>SUB_BOS(614), OKO=>SUB_OKOS(614), D=>SUB_DS(614), SO=>SUB_SOS(614));
	DIV615: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(582), SI=>SUB_SOS(583), BI=>SUB_BOS(614), OKI=>SUB_OKOS(616), BO=>SUB_BOS(615), OKO=>SUB_OKOS(615), D=>SUB_DS(615), SO=>SUB_SOS(615));
	DIV616: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(583), SI=>SUB_SOS(584), BI=>SUB_BOS(615), OKI=>SUB_OKOS(617), BO=>SUB_BOS(616), OKO=>SUB_OKOS(616), D=>SUB_DS(616), SO=>SUB_SOS(616));
	DIV617: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(584), SI=>SUB_SOS(585), BI=>SUB_BOS(616), OKI=>SUB_OKOS(618), BO=>SUB_BOS(617), OKO=>SUB_OKOS(617), D=>SUB_DS(617), SO=>SUB_SOS(617));
	DIV618: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(585), SI=>SUB_SOS(586), BI=>SUB_BOS(617), OKI=>SUB_OKOS(619), BO=>SUB_BOS(618), OKO=>SUB_OKOS(618), D=>SUB_DS(618), SO=>SUB_SOS(618));
	DIV619: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(586), SI=>SUB_SOS(587), BI=>SUB_BOS(618), OKI=>SUB_OKOS(620), BO=>SUB_BOS(619), OKO=>SUB_OKOS(619), D=>SUB_DS(619), SO=>SUB_SOS(619));
	DIV620: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(587), SI=>SUB_SOS(588), BI=>SUB_BOS(619), OKI=>SUB_OKOS(621), BO=>SUB_BOS(620), OKO=>SUB_OKOS(620), D=>SUB_DS(620), SO=>SUB_SOS(620));
	DIV621: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(588), SI=>SUB_SOS(589), BI=>SUB_BOS(620), OKI=>SUB_OKOS(622), BO=>SUB_BOS(621), OKO=>SUB_OKOS(621), D=>SUB_DS(621), SO=>SUB_SOS(621));
	DIV622: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(589), SI=>SUB_SOS(590), BI=>SUB_BOS(621), OKI=>SUB_OKOS(623), BO=>SUB_BOS(622), OKO=>SUB_OKOS(622), D=>SUB_DS(622), SO=>SUB_SOS(622));
	DIV623: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(590), SI=>SUB_SOS(591), BI=>SUB_BOS(622), OKI=>SUB_OKOS(624), BO=>SUB_BOS(623), OKO=>SUB_OKOS(623), D=>SUB_DS(623), SO=>SUB_SOS(623));
	DIV624: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(591), SI=>SUB_SOS(592), BI=>SUB_BOS(623), OKI=>SUB_OKOS(625), BO=>SUB_BOS(624), OKO=>SUB_OKOS(624), D=>SUB_DS(624), SO=>SUB_SOS(624));
	DIV625: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(592), SI=>SUB_SOS(593), BI=>SUB_BOS(624), OKI=>SUB_OKOS(626), BO=>SUB_BOS(625), OKO=>SUB_OKOS(625), D=>SUB_DS(625), SO=>SUB_SOS(625));
	DIV626: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(593), SI=>SUB_SOS(594), BI=>SUB_BOS(625), OKI=>SUB_OKOS(627), BO=>SUB_BOS(626), OKO=>SUB_OKOS(626), D=>SUB_DS(626), SO=>SUB_SOS(626));
	DIV627: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(594), SI=>SUB_SOS(595), BI=>SUB_BOS(626), OKI=>SUB_OKOS(628), BO=>SUB_BOS(627), OKO=>SUB_OKOS(627), D=>SUB_DS(627), SO=>SUB_SOS(627));
	DIV628: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(595), SI=>SUB_SOS(596), BI=>SUB_BOS(627), OKI=>SUB_OKOS(629), BO=>SUB_BOS(628), OKO=>SUB_OKOS(628), D=>SUB_DS(628), SO=>SUB_SOS(628));
	DIV629: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(596), SI=>SUB_SOS(597), BI=>SUB_BOS(628), OKI=>SUB_OKOS(630), BO=>SUB_BOS(629), OKO=>SUB_OKOS(629), D=>SUB_DS(629), SO=>SUB_SOS(629));
	DIV630: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(597), SI=>SUB_SOS(598), BI=>SUB_BOS(629), OKI=>SUB_OKOS(631), BO=>SUB_BOS(630), OKO=>SUB_OKOS(630), D=>SUB_DS(630), SO=>SUB_SOS(630));
	DIV631: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(598), SI=>SUB_SOS(599), BI=>SUB_BOS(630), OKI=>SUB_OKOS(632), BO=>SUB_BOS(631), OKO=>SUB_OKOS(631), D=>SUB_DS(631), SO=>SUB_SOS(631));
	DIV632: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(599), SI=>SUB_SOS(600), BI=>SUB_BOS(631), OKI=>SUB_OKOS(633), BO=>SUB_BOS(632), OKO=>SUB_OKOS(632), D=>SUB_DS(632), SO=>SUB_SOS(632));
	DIV633: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(600), SI=>SUB_SOS(601), BI=>SUB_BOS(632), OKI=>SUB_OKOS(634), BO=>SUB_BOS(633), OKO=>SUB_OKOS(633), D=>SUB_DS(633), SO=>SUB_SOS(633));
	DIV634: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(601), SI=>SUB_SOS(602), BI=>SUB_BOS(633), OKI=>SUB_OKOS(635), BO=>SUB_BOS(634), OKO=>SUB_OKOS(634), D=>SUB_DS(634), SO=>SUB_SOS(634));
	DIV635: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(602), SI=>SUB_SOS(603), BI=>SUB_BOS(634), OKI=>SUB_OKOS(636), BO=>SUB_BOS(635), OKO=>SUB_OKOS(635), D=>SUB_DS(635), SO=>SUB_SOS(635));
	DIV636: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(603), SI=>SUB_SOS(604), BI=>SUB_BOS(635), OKI=>SUB_OKOS(637), BO=>SUB_BOS(636), OKO=>SUB_OKOS(636), D=>SUB_DS(636), SO=>SUB_SOS(636));
	DIV637: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(604), SI=>SUB_SOS(605), BI=>SUB_BOS(636), OKI=>SUB_OKOS(638), BO=>SUB_BOS(637), OKO=>SUB_OKOS(637), D=>SUB_DS(637), SO=>SUB_SOS(637));
	DIV638: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(605), SI=>SUB_SOS(606), BI=>SUB_BOS(637), OKI=>SUB_OKOS(639), BO=>SUB_BOS(638), OKO=>SUB_OKOS(638), D=>SUB_DS(638), SO=>SUB_SOS(638));
	DIV639: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(606), SI=>SUB_SOS(607), BI=>SUB_BOS(638), OKI=>BONS(19), BO=>SUB_BOS(639), OKO=>SUB_OKOS(639), D=>SUB_DS(639), SO=>SUB_SOS(639));

	DIV640: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(11), SI=>SUB_SOS(608), BI=>'0', OKI=>SUB_OKOS(641), BO=>SUB_BOS(640), OKO=>SUB_OKOS(640), D=>SUB_DS(640), SO=>SUB_SOS(640));
	DIV641: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(608), SI=>SUB_SOS(609), BI=>SUB_BOS(640), OKI=>SUB_OKOS(642), BO=>SUB_BOS(641), OKO=>SUB_OKOS(641), D=>SUB_DS(641), SO=>SUB_SOS(641));
	DIV642: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(609), SI=>SUB_SOS(610), BI=>SUB_BOS(641), OKI=>SUB_OKOS(643), BO=>SUB_BOS(642), OKO=>SUB_OKOS(642), D=>SUB_DS(642), SO=>SUB_SOS(642));
	DIV643: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(610), SI=>SUB_SOS(611), BI=>SUB_BOS(642), OKI=>SUB_OKOS(644), BO=>SUB_BOS(643), OKO=>SUB_OKOS(643), D=>SUB_DS(643), SO=>SUB_SOS(643));
	DIV644: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(611), SI=>SUB_SOS(612), BI=>SUB_BOS(643), OKI=>SUB_OKOS(645), BO=>SUB_BOS(644), OKO=>SUB_OKOS(644), D=>SUB_DS(644), SO=>SUB_SOS(644));
	DIV645: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(612), SI=>SUB_SOS(613), BI=>SUB_BOS(644), OKI=>SUB_OKOS(646), BO=>SUB_BOS(645), OKO=>SUB_OKOS(645), D=>SUB_DS(645), SO=>SUB_SOS(645));
	DIV646: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(613), SI=>SUB_SOS(614), BI=>SUB_BOS(645), OKI=>SUB_OKOS(647), BO=>SUB_BOS(646), OKO=>SUB_OKOS(646), D=>SUB_DS(646), SO=>SUB_SOS(646));
	DIV647: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(614), SI=>SUB_SOS(615), BI=>SUB_BOS(646), OKI=>SUB_OKOS(648), BO=>SUB_BOS(647), OKO=>SUB_OKOS(647), D=>SUB_DS(647), SO=>SUB_SOS(647));
	DIV648: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(615), SI=>SUB_SOS(616), BI=>SUB_BOS(647), OKI=>SUB_OKOS(649), BO=>SUB_BOS(648), OKO=>SUB_OKOS(648), D=>SUB_DS(648), SO=>SUB_SOS(648));
	DIV649: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(616), SI=>SUB_SOS(617), BI=>SUB_BOS(648), OKI=>SUB_OKOS(650), BO=>SUB_BOS(649), OKO=>SUB_OKOS(649), D=>SUB_DS(649), SO=>SUB_SOS(649));
	DIV650: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(617), SI=>SUB_SOS(618), BI=>SUB_BOS(649), OKI=>SUB_OKOS(651), BO=>SUB_BOS(650), OKO=>SUB_OKOS(650), D=>SUB_DS(650), SO=>SUB_SOS(650));
	DIV651: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(618), SI=>SUB_SOS(619), BI=>SUB_BOS(650), OKI=>SUB_OKOS(652), BO=>SUB_BOS(651), OKO=>SUB_OKOS(651), D=>SUB_DS(651), SO=>SUB_SOS(651));
	DIV652: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(619), SI=>SUB_SOS(620), BI=>SUB_BOS(651), OKI=>SUB_OKOS(653), BO=>SUB_BOS(652), OKO=>SUB_OKOS(652), D=>SUB_DS(652), SO=>SUB_SOS(652));
	DIV653: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(620), SI=>SUB_SOS(621), BI=>SUB_BOS(652), OKI=>SUB_OKOS(654), BO=>SUB_BOS(653), OKO=>SUB_OKOS(653), D=>SUB_DS(653), SO=>SUB_SOS(653));
	DIV654: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(621), SI=>SUB_SOS(622), BI=>SUB_BOS(653), OKI=>SUB_OKOS(655), BO=>SUB_BOS(654), OKO=>SUB_OKOS(654), D=>SUB_DS(654), SO=>SUB_SOS(654));
	DIV655: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(622), SI=>SUB_SOS(623), BI=>SUB_BOS(654), OKI=>SUB_OKOS(656), BO=>SUB_BOS(655), OKO=>SUB_OKOS(655), D=>SUB_DS(655), SO=>SUB_SOS(655));
	DIV656: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(623), SI=>SUB_SOS(624), BI=>SUB_BOS(655), OKI=>SUB_OKOS(657), BO=>SUB_BOS(656), OKO=>SUB_OKOS(656), D=>SUB_DS(656), SO=>SUB_SOS(656));
	DIV657: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(624), SI=>SUB_SOS(625), BI=>SUB_BOS(656), OKI=>SUB_OKOS(658), BO=>SUB_BOS(657), OKO=>SUB_OKOS(657), D=>SUB_DS(657), SO=>SUB_SOS(657));
	DIV658: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(625), SI=>SUB_SOS(626), BI=>SUB_BOS(657), OKI=>SUB_OKOS(659), BO=>SUB_BOS(658), OKO=>SUB_OKOS(658), D=>SUB_DS(658), SO=>SUB_SOS(658));
	DIV659: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(626), SI=>SUB_SOS(627), BI=>SUB_BOS(658), OKI=>SUB_OKOS(660), BO=>SUB_BOS(659), OKO=>SUB_OKOS(659), D=>SUB_DS(659), SO=>SUB_SOS(659));
	DIV660: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(627), SI=>SUB_SOS(628), BI=>SUB_BOS(659), OKI=>SUB_OKOS(661), BO=>SUB_BOS(660), OKO=>SUB_OKOS(660), D=>SUB_DS(660), SO=>SUB_SOS(660));
	DIV661: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(628), SI=>SUB_SOS(629), BI=>SUB_BOS(660), OKI=>SUB_OKOS(662), BO=>SUB_BOS(661), OKO=>SUB_OKOS(661), D=>SUB_DS(661), SO=>SUB_SOS(661));
	DIV662: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(629), SI=>SUB_SOS(630), BI=>SUB_BOS(661), OKI=>SUB_OKOS(663), BO=>SUB_BOS(662), OKO=>SUB_OKOS(662), D=>SUB_DS(662), SO=>SUB_SOS(662));
	DIV663: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(630), SI=>SUB_SOS(631), BI=>SUB_BOS(662), OKI=>SUB_OKOS(664), BO=>SUB_BOS(663), OKO=>SUB_OKOS(663), D=>SUB_DS(663), SO=>SUB_SOS(663));
	DIV664: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(631), SI=>SUB_SOS(632), BI=>SUB_BOS(663), OKI=>SUB_OKOS(665), BO=>SUB_BOS(664), OKO=>SUB_OKOS(664), D=>SUB_DS(664), SO=>SUB_SOS(664));
	DIV665: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(632), SI=>SUB_SOS(633), BI=>SUB_BOS(664), OKI=>SUB_OKOS(666), BO=>SUB_BOS(665), OKO=>SUB_OKOS(665), D=>SUB_DS(665), SO=>SUB_SOS(665));
	DIV666: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(633), SI=>SUB_SOS(634), BI=>SUB_BOS(665), OKI=>SUB_OKOS(667), BO=>SUB_BOS(666), OKO=>SUB_OKOS(666), D=>SUB_DS(666), SO=>SUB_SOS(666));
	DIV667: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(634), SI=>SUB_SOS(635), BI=>SUB_BOS(666), OKI=>SUB_OKOS(668), BO=>SUB_BOS(667), OKO=>SUB_OKOS(667), D=>SUB_DS(667), SO=>SUB_SOS(667));
	DIV668: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(635), SI=>SUB_SOS(636), BI=>SUB_BOS(667), OKI=>SUB_OKOS(669), BO=>SUB_BOS(668), OKO=>SUB_OKOS(668), D=>SUB_DS(668), SO=>SUB_SOS(668));
	DIV669: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(636), SI=>SUB_SOS(637), BI=>SUB_BOS(668), OKI=>SUB_OKOS(670), BO=>SUB_BOS(669), OKO=>SUB_OKOS(669), D=>SUB_DS(669), SO=>SUB_SOS(669));
	DIV670: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(637), SI=>SUB_SOS(638), BI=>SUB_BOS(669), OKI=>SUB_OKOS(671), BO=>SUB_BOS(670), OKO=>SUB_OKOS(670), D=>SUB_DS(670), SO=>SUB_SOS(670));
	DIV671: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(638), SI=>SUB_SOS(639), BI=>SUB_BOS(670), OKI=>BONS(20), BO=>SUB_BOS(671), OKO=>SUB_OKOS(671), D=>SUB_DS(671), SO=>SUB_SOS(671));

	DIV672: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(10), SI=>SUB_SOS(640), BI=>'0', OKI=>SUB_OKOS(673), BO=>SUB_BOS(672), OKO=>SUB_OKOS(672), D=>SUB_DS(672), SO=>SUB_SOS(672));
	DIV673: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(640), SI=>SUB_SOS(641), BI=>SUB_BOS(672), OKI=>SUB_OKOS(674), BO=>SUB_BOS(673), OKO=>SUB_OKOS(673), D=>SUB_DS(673), SO=>SUB_SOS(673));
	DIV674: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(641), SI=>SUB_SOS(642), BI=>SUB_BOS(673), OKI=>SUB_OKOS(675), BO=>SUB_BOS(674), OKO=>SUB_OKOS(674), D=>SUB_DS(674), SO=>SUB_SOS(674));
	DIV675: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(642), SI=>SUB_SOS(643), BI=>SUB_BOS(674), OKI=>SUB_OKOS(676), BO=>SUB_BOS(675), OKO=>SUB_OKOS(675), D=>SUB_DS(675), SO=>SUB_SOS(675));
	DIV676: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(643), SI=>SUB_SOS(644), BI=>SUB_BOS(675), OKI=>SUB_OKOS(677), BO=>SUB_BOS(676), OKO=>SUB_OKOS(676), D=>SUB_DS(676), SO=>SUB_SOS(676));
	DIV677: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(644), SI=>SUB_SOS(645), BI=>SUB_BOS(676), OKI=>SUB_OKOS(678), BO=>SUB_BOS(677), OKO=>SUB_OKOS(677), D=>SUB_DS(677), SO=>SUB_SOS(677));
	DIV678: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(645), SI=>SUB_SOS(646), BI=>SUB_BOS(677), OKI=>SUB_OKOS(679), BO=>SUB_BOS(678), OKO=>SUB_OKOS(678), D=>SUB_DS(678), SO=>SUB_SOS(678));
	DIV679: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(646), SI=>SUB_SOS(647), BI=>SUB_BOS(678), OKI=>SUB_OKOS(680), BO=>SUB_BOS(679), OKO=>SUB_OKOS(679), D=>SUB_DS(679), SO=>SUB_SOS(679));
	DIV680: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(647), SI=>SUB_SOS(648), BI=>SUB_BOS(679), OKI=>SUB_OKOS(681), BO=>SUB_BOS(680), OKO=>SUB_OKOS(680), D=>SUB_DS(680), SO=>SUB_SOS(680));
	DIV681: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(648), SI=>SUB_SOS(649), BI=>SUB_BOS(680), OKI=>SUB_OKOS(682), BO=>SUB_BOS(681), OKO=>SUB_OKOS(681), D=>SUB_DS(681), SO=>SUB_SOS(681));
	DIV682: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(649), SI=>SUB_SOS(650), BI=>SUB_BOS(681), OKI=>SUB_OKOS(683), BO=>SUB_BOS(682), OKO=>SUB_OKOS(682), D=>SUB_DS(682), SO=>SUB_SOS(682));
	DIV683: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(650), SI=>SUB_SOS(651), BI=>SUB_BOS(682), OKI=>SUB_OKOS(684), BO=>SUB_BOS(683), OKO=>SUB_OKOS(683), D=>SUB_DS(683), SO=>SUB_SOS(683));
	DIV684: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(651), SI=>SUB_SOS(652), BI=>SUB_BOS(683), OKI=>SUB_OKOS(685), BO=>SUB_BOS(684), OKO=>SUB_OKOS(684), D=>SUB_DS(684), SO=>SUB_SOS(684));
	DIV685: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(652), SI=>SUB_SOS(653), BI=>SUB_BOS(684), OKI=>SUB_OKOS(686), BO=>SUB_BOS(685), OKO=>SUB_OKOS(685), D=>SUB_DS(685), SO=>SUB_SOS(685));
	DIV686: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(653), SI=>SUB_SOS(654), BI=>SUB_BOS(685), OKI=>SUB_OKOS(687), BO=>SUB_BOS(686), OKO=>SUB_OKOS(686), D=>SUB_DS(686), SO=>SUB_SOS(686));
	DIV687: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(654), SI=>SUB_SOS(655), BI=>SUB_BOS(686), OKI=>SUB_OKOS(688), BO=>SUB_BOS(687), OKO=>SUB_OKOS(687), D=>SUB_DS(687), SO=>SUB_SOS(687));
	DIV688: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(655), SI=>SUB_SOS(656), BI=>SUB_BOS(687), OKI=>SUB_OKOS(689), BO=>SUB_BOS(688), OKO=>SUB_OKOS(688), D=>SUB_DS(688), SO=>SUB_SOS(688));
	DIV689: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(656), SI=>SUB_SOS(657), BI=>SUB_BOS(688), OKI=>SUB_OKOS(690), BO=>SUB_BOS(689), OKO=>SUB_OKOS(689), D=>SUB_DS(689), SO=>SUB_SOS(689));
	DIV690: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(657), SI=>SUB_SOS(658), BI=>SUB_BOS(689), OKI=>SUB_OKOS(691), BO=>SUB_BOS(690), OKO=>SUB_OKOS(690), D=>SUB_DS(690), SO=>SUB_SOS(690));
	DIV691: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(658), SI=>SUB_SOS(659), BI=>SUB_BOS(690), OKI=>SUB_OKOS(692), BO=>SUB_BOS(691), OKO=>SUB_OKOS(691), D=>SUB_DS(691), SO=>SUB_SOS(691));
	DIV692: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(659), SI=>SUB_SOS(660), BI=>SUB_BOS(691), OKI=>SUB_OKOS(693), BO=>SUB_BOS(692), OKO=>SUB_OKOS(692), D=>SUB_DS(692), SO=>SUB_SOS(692));
	DIV693: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(660), SI=>SUB_SOS(661), BI=>SUB_BOS(692), OKI=>SUB_OKOS(694), BO=>SUB_BOS(693), OKO=>SUB_OKOS(693), D=>SUB_DS(693), SO=>SUB_SOS(693));
	DIV694: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(661), SI=>SUB_SOS(662), BI=>SUB_BOS(693), OKI=>SUB_OKOS(695), BO=>SUB_BOS(694), OKO=>SUB_OKOS(694), D=>SUB_DS(694), SO=>SUB_SOS(694));
	DIV695: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(662), SI=>SUB_SOS(663), BI=>SUB_BOS(694), OKI=>SUB_OKOS(696), BO=>SUB_BOS(695), OKO=>SUB_OKOS(695), D=>SUB_DS(695), SO=>SUB_SOS(695));
	DIV696: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(663), SI=>SUB_SOS(664), BI=>SUB_BOS(695), OKI=>SUB_OKOS(697), BO=>SUB_BOS(696), OKO=>SUB_OKOS(696), D=>SUB_DS(696), SO=>SUB_SOS(696));
	DIV697: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(664), SI=>SUB_SOS(665), BI=>SUB_BOS(696), OKI=>SUB_OKOS(698), BO=>SUB_BOS(697), OKO=>SUB_OKOS(697), D=>SUB_DS(697), SO=>SUB_SOS(697));
	DIV698: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(665), SI=>SUB_SOS(666), BI=>SUB_BOS(697), OKI=>SUB_OKOS(699), BO=>SUB_BOS(698), OKO=>SUB_OKOS(698), D=>SUB_DS(698), SO=>SUB_SOS(698));
	DIV699: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(666), SI=>SUB_SOS(667), BI=>SUB_BOS(698), OKI=>SUB_OKOS(700), BO=>SUB_BOS(699), OKO=>SUB_OKOS(699), D=>SUB_DS(699), SO=>SUB_SOS(699));
	DIV700: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(667), SI=>SUB_SOS(668), BI=>SUB_BOS(699), OKI=>SUB_OKOS(701), BO=>SUB_BOS(700), OKO=>SUB_OKOS(700), D=>SUB_DS(700), SO=>SUB_SOS(700));
	DIV701: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(668), SI=>SUB_SOS(669), BI=>SUB_BOS(700), OKI=>SUB_OKOS(702), BO=>SUB_BOS(701), OKO=>SUB_OKOS(701), D=>SUB_DS(701), SO=>SUB_SOS(701));
	DIV702: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(669), SI=>SUB_SOS(670), BI=>SUB_BOS(701), OKI=>SUB_OKOS(703), BO=>SUB_BOS(702), OKO=>SUB_OKOS(702), D=>SUB_DS(702), SO=>SUB_SOS(702));
	DIV703: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(670), SI=>SUB_SOS(671), BI=>SUB_BOS(702), OKI=>BONS(21), BO=>SUB_BOS(703), OKO=>SUB_OKOS(703), D=>SUB_DS(703), SO=>SUB_SOS(703));

	DIV704: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(9), SI=>SUB_SOS(672), BI=>'0', OKI=>SUB_OKOS(705), BO=>SUB_BOS(704), OKO=>SUB_OKOS(704), D=>SUB_DS(704), SO=>SUB_SOS(704));
	DIV705: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(672), SI=>SUB_SOS(673), BI=>SUB_BOS(704), OKI=>SUB_OKOS(706), BO=>SUB_BOS(705), OKO=>SUB_OKOS(705), D=>SUB_DS(705), SO=>SUB_SOS(705));
	DIV706: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(673), SI=>SUB_SOS(674), BI=>SUB_BOS(705), OKI=>SUB_OKOS(707), BO=>SUB_BOS(706), OKO=>SUB_OKOS(706), D=>SUB_DS(706), SO=>SUB_SOS(706));
	DIV707: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(674), SI=>SUB_SOS(675), BI=>SUB_BOS(706), OKI=>SUB_OKOS(708), BO=>SUB_BOS(707), OKO=>SUB_OKOS(707), D=>SUB_DS(707), SO=>SUB_SOS(707));
	DIV708: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(675), SI=>SUB_SOS(676), BI=>SUB_BOS(707), OKI=>SUB_OKOS(709), BO=>SUB_BOS(708), OKO=>SUB_OKOS(708), D=>SUB_DS(708), SO=>SUB_SOS(708));
	DIV709: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(676), SI=>SUB_SOS(677), BI=>SUB_BOS(708), OKI=>SUB_OKOS(710), BO=>SUB_BOS(709), OKO=>SUB_OKOS(709), D=>SUB_DS(709), SO=>SUB_SOS(709));
	DIV710: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(677), SI=>SUB_SOS(678), BI=>SUB_BOS(709), OKI=>SUB_OKOS(711), BO=>SUB_BOS(710), OKO=>SUB_OKOS(710), D=>SUB_DS(710), SO=>SUB_SOS(710));
	DIV711: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(678), SI=>SUB_SOS(679), BI=>SUB_BOS(710), OKI=>SUB_OKOS(712), BO=>SUB_BOS(711), OKO=>SUB_OKOS(711), D=>SUB_DS(711), SO=>SUB_SOS(711));
	DIV712: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(679), SI=>SUB_SOS(680), BI=>SUB_BOS(711), OKI=>SUB_OKOS(713), BO=>SUB_BOS(712), OKO=>SUB_OKOS(712), D=>SUB_DS(712), SO=>SUB_SOS(712));
	DIV713: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(680), SI=>SUB_SOS(681), BI=>SUB_BOS(712), OKI=>SUB_OKOS(714), BO=>SUB_BOS(713), OKO=>SUB_OKOS(713), D=>SUB_DS(713), SO=>SUB_SOS(713));
	DIV714: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(681), SI=>SUB_SOS(682), BI=>SUB_BOS(713), OKI=>SUB_OKOS(715), BO=>SUB_BOS(714), OKO=>SUB_OKOS(714), D=>SUB_DS(714), SO=>SUB_SOS(714));
	DIV715: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(682), SI=>SUB_SOS(683), BI=>SUB_BOS(714), OKI=>SUB_OKOS(716), BO=>SUB_BOS(715), OKO=>SUB_OKOS(715), D=>SUB_DS(715), SO=>SUB_SOS(715));
	DIV716: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(683), SI=>SUB_SOS(684), BI=>SUB_BOS(715), OKI=>SUB_OKOS(717), BO=>SUB_BOS(716), OKO=>SUB_OKOS(716), D=>SUB_DS(716), SO=>SUB_SOS(716));
	DIV717: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(684), SI=>SUB_SOS(685), BI=>SUB_BOS(716), OKI=>SUB_OKOS(718), BO=>SUB_BOS(717), OKO=>SUB_OKOS(717), D=>SUB_DS(717), SO=>SUB_SOS(717));
	DIV718: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(685), SI=>SUB_SOS(686), BI=>SUB_BOS(717), OKI=>SUB_OKOS(719), BO=>SUB_BOS(718), OKO=>SUB_OKOS(718), D=>SUB_DS(718), SO=>SUB_SOS(718));
	DIV719: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(686), SI=>SUB_SOS(687), BI=>SUB_BOS(718), OKI=>SUB_OKOS(720), BO=>SUB_BOS(719), OKO=>SUB_OKOS(719), D=>SUB_DS(719), SO=>SUB_SOS(719));
	DIV720: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(687), SI=>SUB_SOS(688), BI=>SUB_BOS(719), OKI=>SUB_OKOS(721), BO=>SUB_BOS(720), OKO=>SUB_OKOS(720), D=>SUB_DS(720), SO=>SUB_SOS(720));
	DIV721: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(688), SI=>SUB_SOS(689), BI=>SUB_BOS(720), OKI=>SUB_OKOS(722), BO=>SUB_BOS(721), OKO=>SUB_OKOS(721), D=>SUB_DS(721), SO=>SUB_SOS(721));
	DIV722: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(689), SI=>SUB_SOS(690), BI=>SUB_BOS(721), OKI=>SUB_OKOS(723), BO=>SUB_BOS(722), OKO=>SUB_OKOS(722), D=>SUB_DS(722), SO=>SUB_SOS(722));
	DIV723: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(690), SI=>SUB_SOS(691), BI=>SUB_BOS(722), OKI=>SUB_OKOS(724), BO=>SUB_BOS(723), OKO=>SUB_OKOS(723), D=>SUB_DS(723), SO=>SUB_SOS(723));
	DIV724: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(691), SI=>SUB_SOS(692), BI=>SUB_BOS(723), OKI=>SUB_OKOS(725), BO=>SUB_BOS(724), OKO=>SUB_OKOS(724), D=>SUB_DS(724), SO=>SUB_SOS(724));
	DIV725: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(692), SI=>SUB_SOS(693), BI=>SUB_BOS(724), OKI=>SUB_OKOS(726), BO=>SUB_BOS(725), OKO=>SUB_OKOS(725), D=>SUB_DS(725), SO=>SUB_SOS(725));
	DIV726: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(693), SI=>SUB_SOS(694), BI=>SUB_BOS(725), OKI=>SUB_OKOS(727), BO=>SUB_BOS(726), OKO=>SUB_OKOS(726), D=>SUB_DS(726), SO=>SUB_SOS(726));
	DIV727: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(694), SI=>SUB_SOS(695), BI=>SUB_BOS(726), OKI=>SUB_OKOS(728), BO=>SUB_BOS(727), OKO=>SUB_OKOS(727), D=>SUB_DS(727), SO=>SUB_SOS(727));
	DIV728: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(695), SI=>SUB_SOS(696), BI=>SUB_BOS(727), OKI=>SUB_OKOS(729), BO=>SUB_BOS(728), OKO=>SUB_OKOS(728), D=>SUB_DS(728), SO=>SUB_SOS(728));
	DIV729: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(696), SI=>SUB_SOS(697), BI=>SUB_BOS(728), OKI=>SUB_OKOS(730), BO=>SUB_BOS(729), OKO=>SUB_OKOS(729), D=>SUB_DS(729), SO=>SUB_SOS(729));
	DIV730: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(697), SI=>SUB_SOS(698), BI=>SUB_BOS(729), OKI=>SUB_OKOS(731), BO=>SUB_BOS(730), OKO=>SUB_OKOS(730), D=>SUB_DS(730), SO=>SUB_SOS(730));
	DIV731: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(698), SI=>SUB_SOS(699), BI=>SUB_BOS(730), OKI=>SUB_OKOS(732), BO=>SUB_BOS(731), OKO=>SUB_OKOS(731), D=>SUB_DS(731), SO=>SUB_SOS(731));
	DIV732: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(699), SI=>SUB_SOS(700), BI=>SUB_BOS(731), OKI=>SUB_OKOS(733), BO=>SUB_BOS(732), OKO=>SUB_OKOS(732), D=>SUB_DS(732), SO=>SUB_SOS(732));
	DIV733: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(700), SI=>SUB_SOS(701), BI=>SUB_BOS(732), OKI=>SUB_OKOS(734), BO=>SUB_BOS(733), OKO=>SUB_OKOS(733), D=>SUB_DS(733), SO=>SUB_SOS(733));
	DIV734: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(701), SI=>SUB_SOS(702), BI=>SUB_BOS(733), OKI=>SUB_OKOS(735), BO=>SUB_BOS(734), OKO=>SUB_OKOS(734), D=>SUB_DS(734), SO=>SUB_SOS(734));
	DIV735: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(702), SI=>SUB_SOS(703), BI=>SUB_BOS(734), OKI=>BONS(22), BO=>SUB_BOS(735), OKO=>SUB_OKOS(735), D=>SUB_DS(735), SO=>SUB_SOS(735));

	DIV736: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(8), SI=>SUB_SOS(704), BI=>'0', OKI=>SUB_OKOS(737), BO=>SUB_BOS(736), OKO=>SUB_OKOS(736), D=>SUB_DS(736), SO=>SUB_SOS(736));
	DIV737: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(704), SI=>SUB_SOS(705), BI=>SUB_BOS(736), OKI=>SUB_OKOS(738), BO=>SUB_BOS(737), OKO=>SUB_OKOS(737), D=>SUB_DS(737), SO=>SUB_SOS(737));
	DIV738: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(705), SI=>SUB_SOS(706), BI=>SUB_BOS(737), OKI=>SUB_OKOS(739), BO=>SUB_BOS(738), OKO=>SUB_OKOS(738), D=>SUB_DS(738), SO=>SUB_SOS(738));
	DIV739: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(706), SI=>SUB_SOS(707), BI=>SUB_BOS(738), OKI=>SUB_OKOS(740), BO=>SUB_BOS(739), OKO=>SUB_OKOS(739), D=>SUB_DS(739), SO=>SUB_SOS(739));
	DIV740: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(707), SI=>SUB_SOS(708), BI=>SUB_BOS(739), OKI=>SUB_OKOS(741), BO=>SUB_BOS(740), OKO=>SUB_OKOS(740), D=>SUB_DS(740), SO=>SUB_SOS(740));
	DIV741: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(708), SI=>SUB_SOS(709), BI=>SUB_BOS(740), OKI=>SUB_OKOS(742), BO=>SUB_BOS(741), OKO=>SUB_OKOS(741), D=>SUB_DS(741), SO=>SUB_SOS(741));
	DIV742: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(709), SI=>SUB_SOS(710), BI=>SUB_BOS(741), OKI=>SUB_OKOS(743), BO=>SUB_BOS(742), OKO=>SUB_OKOS(742), D=>SUB_DS(742), SO=>SUB_SOS(742));
	DIV743: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(710), SI=>SUB_SOS(711), BI=>SUB_BOS(742), OKI=>SUB_OKOS(744), BO=>SUB_BOS(743), OKO=>SUB_OKOS(743), D=>SUB_DS(743), SO=>SUB_SOS(743));
	DIV744: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(711), SI=>SUB_SOS(712), BI=>SUB_BOS(743), OKI=>SUB_OKOS(745), BO=>SUB_BOS(744), OKO=>SUB_OKOS(744), D=>SUB_DS(744), SO=>SUB_SOS(744));
	DIV745: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(712), SI=>SUB_SOS(713), BI=>SUB_BOS(744), OKI=>SUB_OKOS(746), BO=>SUB_BOS(745), OKO=>SUB_OKOS(745), D=>SUB_DS(745), SO=>SUB_SOS(745));
	DIV746: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(713), SI=>SUB_SOS(714), BI=>SUB_BOS(745), OKI=>SUB_OKOS(747), BO=>SUB_BOS(746), OKO=>SUB_OKOS(746), D=>SUB_DS(746), SO=>SUB_SOS(746));
	DIV747: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(714), SI=>SUB_SOS(715), BI=>SUB_BOS(746), OKI=>SUB_OKOS(748), BO=>SUB_BOS(747), OKO=>SUB_OKOS(747), D=>SUB_DS(747), SO=>SUB_SOS(747));
	DIV748: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(715), SI=>SUB_SOS(716), BI=>SUB_BOS(747), OKI=>SUB_OKOS(749), BO=>SUB_BOS(748), OKO=>SUB_OKOS(748), D=>SUB_DS(748), SO=>SUB_SOS(748));
	DIV749: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(716), SI=>SUB_SOS(717), BI=>SUB_BOS(748), OKI=>SUB_OKOS(750), BO=>SUB_BOS(749), OKO=>SUB_OKOS(749), D=>SUB_DS(749), SO=>SUB_SOS(749));
	DIV750: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(717), SI=>SUB_SOS(718), BI=>SUB_BOS(749), OKI=>SUB_OKOS(751), BO=>SUB_BOS(750), OKO=>SUB_OKOS(750), D=>SUB_DS(750), SO=>SUB_SOS(750));
	DIV751: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(718), SI=>SUB_SOS(719), BI=>SUB_BOS(750), OKI=>SUB_OKOS(752), BO=>SUB_BOS(751), OKO=>SUB_OKOS(751), D=>SUB_DS(751), SO=>SUB_SOS(751));
	DIV752: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(719), SI=>SUB_SOS(720), BI=>SUB_BOS(751), OKI=>SUB_OKOS(753), BO=>SUB_BOS(752), OKO=>SUB_OKOS(752), D=>SUB_DS(752), SO=>SUB_SOS(752));
	DIV753: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(720), SI=>SUB_SOS(721), BI=>SUB_BOS(752), OKI=>SUB_OKOS(754), BO=>SUB_BOS(753), OKO=>SUB_OKOS(753), D=>SUB_DS(753), SO=>SUB_SOS(753));
	DIV754: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(721), SI=>SUB_SOS(722), BI=>SUB_BOS(753), OKI=>SUB_OKOS(755), BO=>SUB_BOS(754), OKO=>SUB_OKOS(754), D=>SUB_DS(754), SO=>SUB_SOS(754));
	DIV755: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(722), SI=>SUB_SOS(723), BI=>SUB_BOS(754), OKI=>SUB_OKOS(756), BO=>SUB_BOS(755), OKO=>SUB_OKOS(755), D=>SUB_DS(755), SO=>SUB_SOS(755));
	DIV756: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(723), SI=>SUB_SOS(724), BI=>SUB_BOS(755), OKI=>SUB_OKOS(757), BO=>SUB_BOS(756), OKO=>SUB_OKOS(756), D=>SUB_DS(756), SO=>SUB_SOS(756));
	DIV757: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(724), SI=>SUB_SOS(725), BI=>SUB_BOS(756), OKI=>SUB_OKOS(758), BO=>SUB_BOS(757), OKO=>SUB_OKOS(757), D=>SUB_DS(757), SO=>SUB_SOS(757));
	DIV758: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(725), SI=>SUB_SOS(726), BI=>SUB_BOS(757), OKI=>SUB_OKOS(759), BO=>SUB_BOS(758), OKO=>SUB_OKOS(758), D=>SUB_DS(758), SO=>SUB_SOS(758));
	DIV759: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(726), SI=>SUB_SOS(727), BI=>SUB_BOS(758), OKI=>SUB_OKOS(760), BO=>SUB_BOS(759), OKO=>SUB_OKOS(759), D=>SUB_DS(759), SO=>SUB_SOS(759));
	DIV760: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(727), SI=>SUB_SOS(728), BI=>SUB_BOS(759), OKI=>SUB_OKOS(761), BO=>SUB_BOS(760), OKO=>SUB_OKOS(760), D=>SUB_DS(760), SO=>SUB_SOS(760));
	DIV761: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(728), SI=>SUB_SOS(729), BI=>SUB_BOS(760), OKI=>SUB_OKOS(762), BO=>SUB_BOS(761), OKO=>SUB_OKOS(761), D=>SUB_DS(761), SO=>SUB_SOS(761));
	DIV762: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(729), SI=>SUB_SOS(730), BI=>SUB_BOS(761), OKI=>SUB_OKOS(763), BO=>SUB_BOS(762), OKO=>SUB_OKOS(762), D=>SUB_DS(762), SO=>SUB_SOS(762));
	DIV763: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(730), SI=>SUB_SOS(731), BI=>SUB_BOS(762), OKI=>SUB_OKOS(764), BO=>SUB_BOS(763), OKO=>SUB_OKOS(763), D=>SUB_DS(763), SO=>SUB_SOS(763));
	DIV764: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(731), SI=>SUB_SOS(732), BI=>SUB_BOS(763), OKI=>SUB_OKOS(765), BO=>SUB_BOS(764), OKO=>SUB_OKOS(764), D=>SUB_DS(764), SO=>SUB_SOS(764));
	DIV765: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(732), SI=>SUB_SOS(733), BI=>SUB_BOS(764), OKI=>SUB_OKOS(766), BO=>SUB_BOS(765), OKO=>SUB_OKOS(765), D=>SUB_DS(765), SO=>SUB_SOS(765));
	DIV766: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(733), SI=>SUB_SOS(734), BI=>SUB_BOS(765), OKI=>SUB_OKOS(767), BO=>SUB_BOS(766), OKO=>SUB_OKOS(766), D=>SUB_DS(766), SO=>SUB_SOS(766));
	DIV767: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(734), SI=>SUB_SOS(735), BI=>SUB_BOS(766), OKI=>BONS(23), BO=>SUB_BOS(767), OKO=>SUB_OKOS(767), D=>SUB_DS(767), SO=>SUB_SOS(767));

	DIV768: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(7), SI=>SUB_SOS(736), BI=>'0', OKI=>SUB_OKOS(769), BO=>SUB_BOS(768), OKO=>SUB_OKOS(768), D=>SUB_DS(768), SO=>SUB_SOS(768));
	DIV769: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(736), SI=>SUB_SOS(737), BI=>SUB_BOS(768), OKI=>SUB_OKOS(770), BO=>SUB_BOS(769), OKO=>SUB_OKOS(769), D=>SUB_DS(769), SO=>SUB_SOS(769));
	DIV770: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(737), SI=>SUB_SOS(738), BI=>SUB_BOS(769), OKI=>SUB_OKOS(771), BO=>SUB_BOS(770), OKO=>SUB_OKOS(770), D=>SUB_DS(770), SO=>SUB_SOS(770));
	DIV771: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(738), SI=>SUB_SOS(739), BI=>SUB_BOS(770), OKI=>SUB_OKOS(772), BO=>SUB_BOS(771), OKO=>SUB_OKOS(771), D=>SUB_DS(771), SO=>SUB_SOS(771));
	DIV772: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(739), SI=>SUB_SOS(740), BI=>SUB_BOS(771), OKI=>SUB_OKOS(773), BO=>SUB_BOS(772), OKO=>SUB_OKOS(772), D=>SUB_DS(772), SO=>SUB_SOS(772));
	DIV773: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(740), SI=>SUB_SOS(741), BI=>SUB_BOS(772), OKI=>SUB_OKOS(774), BO=>SUB_BOS(773), OKO=>SUB_OKOS(773), D=>SUB_DS(773), SO=>SUB_SOS(773));
	DIV774: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(741), SI=>SUB_SOS(742), BI=>SUB_BOS(773), OKI=>SUB_OKOS(775), BO=>SUB_BOS(774), OKO=>SUB_OKOS(774), D=>SUB_DS(774), SO=>SUB_SOS(774));
	DIV775: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(742), SI=>SUB_SOS(743), BI=>SUB_BOS(774), OKI=>SUB_OKOS(776), BO=>SUB_BOS(775), OKO=>SUB_OKOS(775), D=>SUB_DS(775), SO=>SUB_SOS(775));
	DIV776: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(743), SI=>SUB_SOS(744), BI=>SUB_BOS(775), OKI=>SUB_OKOS(777), BO=>SUB_BOS(776), OKO=>SUB_OKOS(776), D=>SUB_DS(776), SO=>SUB_SOS(776));
	DIV777: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(744), SI=>SUB_SOS(745), BI=>SUB_BOS(776), OKI=>SUB_OKOS(778), BO=>SUB_BOS(777), OKO=>SUB_OKOS(777), D=>SUB_DS(777), SO=>SUB_SOS(777));
	DIV778: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(745), SI=>SUB_SOS(746), BI=>SUB_BOS(777), OKI=>SUB_OKOS(779), BO=>SUB_BOS(778), OKO=>SUB_OKOS(778), D=>SUB_DS(778), SO=>SUB_SOS(778));
	DIV779: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(746), SI=>SUB_SOS(747), BI=>SUB_BOS(778), OKI=>SUB_OKOS(780), BO=>SUB_BOS(779), OKO=>SUB_OKOS(779), D=>SUB_DS(779), SO=>SUB_SOS(779));
	DIV780: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(747), SI=>SUB_SOS(748), BI=>SUB_BOS(779), OKI=>SUB_OKOS(781), BO=>SUB_BOS(780), OKO=>SUB_OKOS(780), D=>SUB_DS(780), SO=>SUB_SOS(780));
	DIV781: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(748), SI=>SUB_SOS(749), BI=>SUB_BOS(780), OKI=>SUB_OKOS(782), BO=>SUB_BOS(781), OKO=>SUB_OKOS(781), D=>SUB_DS(781), SO=>SUB_SOS(781));
	DIV782: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(749), SI=>SUB_SOS(750), BI=>SUB_BOS(781), OKI=>SUB_OKOS(783), BO=>SUB_BOS(782), OKO=>SUB_OKOS(782), D=>SUB_DS(782), SO=>SUB_SOS(782));
	DIV783: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(750), SI=>SUB_SOS(751), BI=>SUB_BOS(782), OKI=>SUB_OKOS(784), BO=>SUB_BOS(783), OKO=>SUB_OKOS(783), D=>SUB_DS(783), SO=>SUB_SOS(783));
	DIV784: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(751), SI=>SUB_SOS(752), BI=>SUB_BOS(783), OKI=>SUB_OKOS(785), BO=>SUB_BOS(784), OKO=>SUB_OKOS(784), D=>SUB_DS(784), SO=>SUB_SOS(784));
	DIV785: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(752), SI=>SUB_SOS(753), BI=>SUB_BOS(784), OKI=>SUB_OKOS(786), BO=>SUB_BOS(785), OKO=>SUB_OKOS(785), D=>SUB_DS(785), SO=>SUB_SOS(785));
	DIV786: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(753), SI=>SUB_SOS(754), BI=>SUB_BOS(785), OKI=>SUB_OKOS(787), BO=>SUB_BOS(786), OKO=>SUB_OKOS(786), D=>SUB_DS(786), SO=>SUB_SOS(786));
	DIV787: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(754), SI=>SUB_SOS(755), BI=>SUB_BOS(786), OKI=>SUB_OKOS(788), BO=>SUB_BOS(787), OKO=>SUB_OKOS(787), D=>SUB_DS(787), SO=>SUB_SOS(787));
	DIV788: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(755), SI=>SUB_SOS(756), BI=>SUB_BOS(787), OKI=>SUB_OKOS(789), BO=>SUB_BOS(788), OKO=>SUB_OKOS(788), D=>SUB_DS(788), SO=>SUB_SOS(788));
	DIV789: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(756), SI=>SUB_SOS(757), BI=>SUB_BOS(788), OKI=>SUB_OKOS(790), BO=>SUB_BOS(789), OKO=>SUB_OKOS(789), D=>SUB_DS(789), SO=>SUB_SOS(789));
	DIV790: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(757), SI=>SUB_SOS(758), BI=>SUB_BOS(789), OKI=>SUB_OKOS(791), BO=>SUB_BOS(790), OKO=>SUB_OKOS(790), D=>SUB_DS(790), SO=>SUB_SOS(790));
	DIV791: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(758), SI=>SUB_SOS(759), BI=>SUB_BOS(790), OKI=>SUB_OKOS(792), BO=>SUB_BOS(791), OKO=>SUB_OKOS(791), D=>SUB_DS(791), SO=>SUB_SOS(791));
	DIV792: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(759), SI=>SUB_SOS(760), BI=>SUB_BOS(791), OKI=>SUB_OKOS(793), BO=>SUB_BOS(792), OKO=>SUB_OKOS(792), D=>SUB_DS(792), SO=>SUB_SOS(792));
	DIV793: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(760), SI=>SUB_SOS(761), BI=>SUB_BOS(792), OKI=>SUB_OKOS(794), BO=>SUB_BOS(793), OKO=>SUB_OKOS(793), D=>SUB_DS(793), SO=>SUB_SOS(793));
	DIV794: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(761), SI=>SUB_SOS(762), BI=>SUB_BOS(793), OKI=>SUB_OKOS(795), BO=>SUB_BOS(794), OKO=>SUB_OKOS(794), D=>SUB_DS(794), SO=>SUB_SOS(794));
	DIV795: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(762), SI=>SUB_SOS(763), BI=>SUB_BOS(794), OKI=>SUB_OKOS(796), BO=>SUB_BOS(795), OKO=>SUB_OKOS(795), D=>SUB_DS(795), SO=>SUB_SOS(795));
	DIV796: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(763), SI=>SUB_SOS(764), BI=>SUB_BOS(795), OKI=>SUB_OKOS(797), BO=>SUB_BOS(796), OKO=>SUB_OKOS(796), D=>SUB_DS(796), SO=>SUB_SOS(796));
	DIV797: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(764), SI=>SUB_SOS(765), BI=>SUB_BOS(796), OKI=>SUB_OKOS(798), BO=>SUB_BOS(797), OKO=>SUB_OKOS(797), D=>SUB_DS(797), SO=>SUB_SOS(797));
	DIV798: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(765), SI=>SUB_SOS(766), BI=>SUB_BOS(797), OKI=>SUB_OKOS(799), BO=>SUB_BOS(798), OKO=>SUB_OKOS(798), D=>SUB_DS(798), SO=>SUB_SOS(798));
	DIV799: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(766), SI=>SUB_SOS(767), BI=>SUB_BOS(798), OKI=>BONS(24), BO=>SUB_BOS(799), OKO=>SUB_OKOS(799), D=>SUB_DS(799), SO=>SUB_SOS(799));

	DIV800: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(6), SI=>SUB_SOS(768), BI=>'0', OKI=>SUB_OKOS(801), BO=>SUB_BOS(800), OKO=>SUB_OKOS(800), D=>SUB_DS(800), SO=>SUB_SOS(800));
	DIV801: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(768), SI=>SUB_SOS(769), BI=>SUB_BOS(800), OKI=>SUB_OKOS(802), BO=>SUB_BOS(801), OKO=>SUB_OKOS(801), D=>SUB_DS(801), SO=>SUB_SOS(801));
	DIV802: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(769), SI=>SUB_SOS(770), BI=>SUB_BOS(801), OKI=>SUB_OKOS(803), BO=>SUB_BOS(802), OKO=>SUB_OKOS(802), D=>SUB_DS(802), SO=>SUB_SOS(802));
	DIV803: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(770), SI=>SUB_SOS(771), BI=>SUB_BOS(802), OKI=>SUB_OKOS(804), BO=>SUB_BOS(803), OKO=>SUB_OKOS(803), D=>SUB_DS(803), SO=>SUB_SOS(803));
	DIV804: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(771), SI=>SUB_SOS(772), BI=>SUB_BOS(803), OKI=>SUB_OKOS(805), BO=>SUB_BOS(804), OKO=>SUB_OKOS(804), D=>SUB_DS(804), SO=>SUB_SOS(804));
	DIV805: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(772), SI=>SUB_SOS(773), BI=>SUB_BOS(804), OKI=>SUB_OKOS(806), BO=>SUB_BOS(805), OKO=>SUB_OKOS(805), D=>SUB_DS(805), SO=>SUB_SOS(805));
	DIV806: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(773), SI=>SUB_SOS(774), BI=>SUB_BOS(805), OKI=>SUB_OKOS(807), BO=>SUB_BOS(806), OKO=>SUB_OKOS(806), D=>SUB_DS(806), SO=>SUB_SOS(806));
	DIV807: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(774), SI=>SUB_SOS(775), BI=>SUB_BOS(806), OKI=>SUB_OKOS(808), BO=>SUB_BOS(807), OKO=>SUB_OKOS(807), D=>SUB_DS(807), SO=>SUB_SOS(807));
	DIV808: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(775), SI=>SUB_SOS(776), BI=>SUB_BOS(807), OKI=>SUB_OKOS(809), BO=>SUB_BOS(808), OKO=>SUB_OKOS(808), D=>SUB_DS(808), SO=>SUB_SOS(808));
	DIV809: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(776), SI=>SUB_SOS(777), BI=>SUB_BOS(808), OKI=>SUB_OKOS(810), BO=>SUB_BOS(809), OKO=>SUB_OKOS(809), D=>SUB_DS(809), SO=>SUB_SOS(809));
	DIV810: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(777), SI=>SUB_SOS(778), BI=>SUB_BOS(809), OKI=>SUB_OKOS(811), BO=>SUB_BOS(810), OKO=>SUB_OKOS(810), D=>SUB_DS(810), SO=>SUB_SOS(810));
	DIV811: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(778), SI=>SUB_SOS(779), BI=>SUB_BOS(810), OKI=>SUB_OKOS(812), BO=>SUB_BOS(811), OKO=>SUB_OKOS(811), D=>SUB_DS(811), SO=>SUB_SOS(811));
	DIV812: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(779), SI=>SUB_SOS(780), BI=>SUB_BOS(811), OKI=>SUB_OKOS(813), BO=>SUB_BOS(812), OKO=>SUB_OKOS(812), D=>SUB_DS(812), SO=>SUB_SOS(812));
	DIV813: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(780), SI=>SUB_SOS(781), BI=>SUB_BOS(812), OKI=>SUB_OKOS(814), BO=>SUB_BOS(813), OKO=>SUB_OKOS(813), D=>SUB_DS(813), SO=>SUB_SOS(813));
	DIV814: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(781), SI=>SUB_SOS(782), BI=>SUB_BOS(813), OKI=>SUB_OKOS(815), BO=>SUB_BOS(814), OKO=>SUB_OKOS(814), D=>SUB_DS(814), SO=>SUB_SOS(814));
	DIV815: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(782), SI=>SUB_SOS(783), BI=>SUB_BOS(814), OKI=>SUB_OKOS(816), BO=>SUB_BOS(815), OKO=>SUB_OKOS(815), D=>SUB_DS(815), SO=>SUB_SOS(815));
	DIV816: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(783), SI=>SUB_SOS(784), BI=>SUB_BOS(815), OKI=>SUB_OKOS(817), BO=>SUB_BOS(816), OKO=>SUB_OKOS(816), D=>SUB_DS(816), SO=>SUB_SOS(816));
	DIV817: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(784), SI=>SUB_SOS(785), BI=>SUB_BOS(816), OKI=>SUB_OKOS(818), BO=>SUB_BOS(817), OKO=>SUB_OKOS(817), D=>SUB_DS(817), SO=>SUB_SOS(817));
	DIV818: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(785), SI=>SUB_SOS(786), BI=>SUB_BOS(817), OKI=>SUB_OKOS(819), BO=>SUB_BOS(818), OKO=>SUB_OKOS(818), D=>SUB_DS(818), SO=>SUB_SOS(818));
	DIV819: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(786), SI=>SUB_SOS(787), BI=>SUB_BOS(818), OKI=>SUB_OKOS(820), BO=>SUB_BOS(819), OKO=>SUB_OKOS(819), D=>SUB_DS(819), SO=>SUB_SOS(819));
	DIV820: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(787), SI=>SUB_SOS(788), BI=>SUB_BOS(819), OKI=>SUB_OKOS(821), BO=>SUB_BOS(820), OKO=>SUB_OKOS(820), D=>SUB_DS(820), SO=>SUB_SOS(820));
	DIV821: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(788), SI=>SUB_SOS(789), BI=>SUB_BOS(820), OKI=>SUB_OKOS(822), BO=>SUB_BOS(821), OKO=>SUB_OKOS(821), D=>SUB_DS(821), SO=>SUB_SOS(821));
	DIV822: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(789), SI=>SUB_SOS(790), BI=>SUB_BOS(821), OKI=>SUB_OKOS(823), BO=>SUB_BOS(822), OKO=>SUB_OKOS(822), D=>SUB_DS(822), SO=>SUB_SOS(822));
	DIV823: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(790), SI=>SUB_SOS(791), BI=>SUB_BOS(822), OKI=>SUB_OKOS(824), BO=>SUB_BOS(823), OKO=>SUB_OKOS(823), D=>SUB_DS(823), SO=>SUB_SOS(823));
	DIV824: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(791), SI=>SUB_SOS(792), BI=>SUB_BOS(823), OKI=>SUB_OKOS(825), BO=>SUB_BOS(824), OKO=>SUB_OKOS(824), D=>SUB_DS(824), SO=>SUB_SOS(824));
	DIV825: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(792), SI=>SUB_SOS(793), BI=>SUB_BOS(824), OKI=>SUB_OKOS(826), BO=>SUB_BOS(825), OKO=>SUB_OKOS(825), D=>SUB_DS(825), SO=>SUB_SOS(825));
	DIV826: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(793), SI=>SUB_SOS(794), BI=>SUB_BOS(825), OKI=>SUB_OKOS(827), BO=>SUB_BOS(826), OKO=>SUB_OKOS(826), D=>SUB_DS(826), SO=>SUB_SOS(826));
	DIV827: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(794), SI=>SUB_SOS(795), BI=>SUB_BOS(826), OKI=>SUB_OKOS(828), BO=>SUB_BOS(827), OKO=>SUB_OKOS(827), D=>SUB_DS(827), SO=>SUB_SOS(827));
	DIV828: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(795), SI=>SUB_SOS(796), BI=>SUB_BOS(827), OKI=>SUB_OKOS(829), BO=>SUB_BOS(828), OKO=>SUB_OKOS(828), D=>SUB_DS(828), SO=>SUB_SOS(828));
	DIV829: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(796), SI=>SUB_SOS(797), BI=>SUB_BOS(828), OKI=>SUB_OKOS(830), BO=>SUB_BOS(829), OKO=>SUB_OKOS(829), D=>SUB_DS(829), SO=>SUB_SOS(829));
	DIV830: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(797), SI=>SUB_SOS(798), BI=>SUB_BOS(829), OKI=>SUB_OKOS(831), BO=>SUB_BOS(830), OKO=>SUB_OKOS(830), D=>SUB_DS(830), SO=>SUB_SOS(830));
	DIV831: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(798), SI=>SUB_SOS(799), BI=>SUB_BOS(830), OKI=>BONS(25), BO=>SUB_BOS(831), OKO=>SUB_OKOS(831), D=>SUB_DS(831), SO=>SUB_SOS(831));

	DIV832: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(5), SI=>SUB_SOS(800), BI=>'0', OKI=>SUB_OKOS(833), BO=>SUB_BOS(832), OKO=>SUB_OKOS(832), D=>SUB_DS(832), SO=>SUB_SOS(832));
	DIV833: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(800), SI=>SUB_SOS(801), BI=>SUB_BOS(832), OKI=>SUB_OKOS(834), BO=>SUB_BOS(833), OKO=>SUB_OKOS(833), D=>SUB_DS(833), SO=>SUB_SOS(833));
	DIV834: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(801), SI=>SUB_SOS(802), BI=>SUB_BOS(833), OKI=>SUB_OKOS(835), BO=>SUB_BOS(834), OKO=>SUB_OKOS(834), D=>SUB_DS(834), SO=>SUB_SOS(834));
	DIV835: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(802), SI=>SUB_SOS(803), BI=>SUB_BOS(834), OKI=>SUB_OKOS(836), BO=>SUB_BOS(835), OKO=>SUB_OKOS(835), D=>SUB_DS(835), SO=>SUB_SOS(835));
	DIV836: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(803), SI=>SUB_SOS(804), BI=>SUB_BOS(835), OKI=>SUB_OKOS(837), BO=>SUB_BOS(836), OKO=>SUB_OKOS(836), D=>SUB_DS(836), SO=>SUB_SOS(836));
	DIV837: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(804), SI=>SUB_SOS(805), BI=>SUB_BOS(836), OKI=>SUB_OKOS(838), BO=>SUB_BOS(837), OKO=>SUB_OKOS(837), D=>SUB_DS(837), SO=>SUB_SOS(837));
	DIV838: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(805), SI=>SUB_SOS(806), BI=>SUB_BOS(837), OKI=>SUB_OKOS(839), BO=>SUB_BOS(838), OKO=>SUB_OKOS(838), D=>SUB_DS(838), SO=>SUB_SOS(838));
	DIV839: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(806), SI=>SUB_SOS(807), BI=>SUB_BOS(838), OKI=>SUB_OKOS(840), BO=>SUB_BOS(839), OKO=>SUB_OKOS(839), D=>SUB_DS(839), SO=>SUB_SOS(839));
	DIV840: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(807), SI=>SUB_SOS(808), BI=>SUB_BOS(839), OKI=>SUB_OKOS(841), BO=>SUB_BOS(840), OKO=>SUB_OKOS(840), D=>SUB_DS(840), SO=>SUB_SOS(840));
	DIV841: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(808), SI=>SUB_SOS(809), BI=>SUB_BOS(840), OKI=>SUB_OKOS(842), BO=>SUB_BOS(841), OKO=>SUB_OKOS(841), D=>SUB_DS(841), SO=>SUB_SOS(841));
	DIV842: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(809), SI=>SUB_SOS(810), BI=>SUB_BOS(841), OKI=>SUB_OKOS(843), BO=>SUB_BOS(842), OKO=>SUB_OKOS(842), D=>SUB_DS(842), SO=>SUB_SOS(842));
	DIV843: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(810), SI=>SUB_SOS(811), BI=>SUB_BOS(842), OKI=>SUB_OKOS(844), BO=>SUB_BOS(843), OKO=>SUB_OKOS(843), D=>SUB_DS(843), SO=>SUB_SOS(843));
	DIV844: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(811), SI=>SUB_SOS(812), BI=>SUB_BOS(843), OKI=>SUB_OKOS(845), BO=>SUB_BOS(844), OKO=>SUB_OKOS(844), D=>SUB_DS(844), SO=>SUB_SOS(844));
	DIV845: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(812), SI=>SUB_SOS(813), BI=>SUB_BOS(844), OKI=>SUB_OKOS(846), BO=>SUB_BOS(845), OKO=>SUB_OKOS(845), D=>SUB_DS(845), SO=>SUB_SOS(845));
	DIV846: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(813), SI=>SUB_SOS(814), BI=>SUB_BOS(845), OKI=>SUB_OKOS(847), BO=>SUB_BOS(846), OKO=>SUB_OKOS(846), D=>SUB_DS(846), SO=>SUB_SOS(846));
	DIV847: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(814), SI=>SUB_SOS(815), BI=>SUB_BOS(846), OKI=>SUB_OKOS(848), BO=>SUB_BOS(847), OKO=>SUB_OKOS(847), D=>SUB_DS(847), SO=>SUB_SOS(847));
	DIV848: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(815), SI=>SUB_SOS(816), BI=>SUB_BOS(847), OKI=>SUB_OKOS(849), BO=>SUB_BOS(848), OKO=>SUB_OKOS(848), D=>SUB_DS(848), SO=>SUB_SOS(848));
	DIV849: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(816), SI=>SUB_SOS(817), BI=>SUB_BOS(848), OKI=>SUB_OKOS(850), BO=>SUB_BOS(849), OKO=>SUB_OKOS(849), D=>SUB_DS(849), SO=>SUB_SOS(849));
	DIV850: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(817), SI=>SUB_SOS(818), BI=>SUB_BOS(849), OKI=>SUB_OKOS(851), BO=>SUB_BOS(850), OKO=>SUB_OKOS(850), D=>SUB_DS(850), SO=>SUB_SOS(850));
	DIV851: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(818), SI=>SUB_SOS(819), BI=>SUB_BOS(850), OKI=>SUB_OKOS(852), BO=>SUB_BOS(851), OKO=>SUB_OKOS(851), D=>SUB_DS(851), SO=>SUB_SOS(851));
	DIV852: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(819), SI=>SUB_SOS(820), BI=>SUB_BOS(851), OKI=>SUB_OKOS(853), BO=>SUB_BOS(852), OKO=>SUB_OKOS(852), D=>SUB_DS(852), SO=>SUB_SOS(852));
	DIV853: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(820), SI=>SUB_SOS(821), BI=>SUB_BOS(852), OKI=>SUB_OKOS(854), BO=>SUB_BOS(853), OKO=>SUB_OKOS(853), D=>SUB_DS(853), SO=>SUB_SOS(853));
	DIV854: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(821), SI=>SUB_SOS(822), BI=>SUB_BOS(853), OKI=>SUB_OKOS(855), BO=>SUB_BOS(854), OKO=>SUB_OKOS(854), D=>SUB_DS(854), SO=>SUB_SOS(854));
	DIV855: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(822), SI=>SUB_SOS(823), BI=>SUB_BOS(854), OKI=>SUB_OKOS(856), BO=>SUB_BOS(855), OKO=>SUB_OKOS(855), D=>SUB_DS(855), SO=>SUB_SOS(855));
	DIV856: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(823), SI=>SUB_SOS(824), BI=>SUB_BOS(855), OKI=>SUB_OKOS(857), BO=>SUB_BOS(856), OKO=>SUB_OKOS(856), D=>SUB_DS(856), SO=>SUB_SOS(856));
	DIV857: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(824), SI=>SUB_SOS(825), BI=>SUB_BOS(856), OKI=>SUB_OKOS(858), BO=>SUB_BOS(857), OKO=>SUB_OKOS(857), D=>SUB_DS(857), SO=>SUB_SOS(857));
	DIV858: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(825), SI=>SUB_SOS(826), BI=>SUB_BOS(857), OKI=>SUB_OKOS(859), BO=>SUB_BOS(858), OKO=>SUB_OKOS(858), D=>SUB_DS(858), SO=>SUB_SOS(858));
	DIV859: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(826), SI=>SUB_SOS(827), BI=>SUB_BOS(858), OKI=>SUB_OKOS(860), BO=>SUB_BOS(859), OKO=>SUB_OKOS(859), D=>SUB_DS(859), SO=>SUB_SOS(859));
	DIV860: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(827), SI=>SUB_SOS(828), BI=>SUB_BOS(859), OKI=>SUB_OKOS(861), BO=>SUB_BOS(860), OKO=>SUB_OKOS(860), D=>SUB_DS(860), SO=>SUB_SOS(860));
	DIV861: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(828), SI=>SUB_SOS(829), BI=>SUB_BOS(860), OKI=>SUB_OKOS(862), BO=>SUB_BOS(861), OKO=>SUB_OKOS(861), D=>SUB_DS(861), SO=>SUB_SOS(861));
	DIV862: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(829), SI=>SUB_SOS(830), BI=>SUB_BOS(861), OKI=>SUB_OKOS(863), BO=>SUB_BOS(862), OKO=>SUB_OKOS(862), D=>SUB_DS(862), SO=>SUB_SOS(862));
	DIV863: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(830), SI=>SUB_SOS(831), BI=>SUB_BOS(862), OKI=>BONS(26), BO=>SUB_BOS(863), OKO=>SUB_OKOS(863), D=>SUB_DS(863), SO=>SUB_SOS(863));

	DIV864: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(4), SI=>SUB_SOS(832), BI=>'0', OKI=>SUB_OKOS(865), BO=>SUB_BOS(864), OKO=>SUB_OKOS(864), D=>SUB_DS(864), SO=>SUB_SOS(864));
	DIV865: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(832), SI=>SUB_SOS(833), BI=>SUB_BOS(864), OKI=>SUB_OKOS(866), BO=>SUB_BOS(865), OKO=>SUB_OKOS(865), D=>SUB_DS(865), SO=>SUB_SOS(865));
	DIV866: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(833), SI=>SUB_SOS(834), BI=>SUB_BOS(865), OKI=>SUB_OKOS(867), BO=>SUB_BOS(866), OKO=>SUB_OKOS(866), D=>SUB_DS(866), SO=>SUB_SOS(866));
	DIV867: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(834), SI=>SUB_SOS(835), BI=>SUB_BOS(866), OKI=>SUB_OKOS(868), BO=>SUB_BOS(867), OKO=>SUB_OKOS(867), D=>SUB_DS(867), SO=>SUB_SOS(867));
	DIV868: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(835), SI=>SUB_SOS(836), BI=>SUB_BOS(867), OKI=>SUB_OKOS(869), BO=>SUB_BOS(868), OKO=>SUB_OKOS(868), D=>SUB_DS(868), SO=>SUB_SOS(868));
	DIV869: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(836), SI=>SUB_SOS(837), BI=>SUB_BOS(868), OKI=>SUB_OKOS(870), BO=>SUB_BOS(869), OKO=>SUB_OKOS(869), D=>SUB_DS(869), SO=>SUB_SOS(869));
	DIV870: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(837), SI=>SUB_SOS(838), BI=>SUB_BOS(869), OKI=>SUB_OKOS(871), BO=>SUB_BOS(870), OKO=>SUB_OKOS(870), D=>SUB_DS(870), SO=>SUB_SOS(870));
	DIV871: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(838), SI=>SUB_SOS(839), BI=>SUB_BOS(870), OKI=>SUB_OKOS(872), BO=>SUB_BOS(871), OKO=>SUB_OKOS(871), D=>SUB_DS(871), SO=>SUB_SOS(871));
	DIV872: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(839), SI=>SUB_SOS(840), BI=>SUB_BOS(871), OKI=>SUB_OKOS(873), BO=>SUB_BOS(872), OKO=>SUB_OKOS(872), D=>SUB_DS(872), SO=>SUB_SOS(872));
	DIV873: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(840), SI=>SUB_SOS(841), BI=>SUB_BOS(872), OKI=>SUB_OKOS(874), BO=>SUB_BOS(873), OKO=>SUB_OKOS(873), D=>SUB_DS(873), SO=>SUB_SOS(873));
	DIV874: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(841), SI=>SUB_SOS(842), BI=>SUB_BOS(873), OKI=>SUB_OKOS(875), BO=>SUB_BOS(874), OKO=>SUB_OKOS(874), D=>SUB_DS(874), SO=>SUB_SOS(874));
	DIV875: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(842), SI=>SUB_SOS(843), BI=>SUB_BOS(874), OKI=>SUB_OKOS(876), BO=>SUB_BOS(875), OKO=>SUB_OKOS(875), D=>SUB_DS(875), SO=>SUB_SOS(875));
	DIV876: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(843), SI=>SUB_SOS(844), BI=>SUB_BOS(875), OKI=>SUB_OKOS(877), BO=>SUB_BOS(876), OKO=>SUB_OKOS(876), D=>SUB_DS(876), SO=>SUB_SOS(876));
	DIV877: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(844), SI=>SUB_SOS(845), BI=>SUB_BOS(876), OKI=>SUB_OKOS(878), BO=>SUB_BOS(877), OKO=>SUB_OKOS(877), D=>SUB_DS(877), SO=>SUB_SOS(877));
	DIV878: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(845), SI=>SUB_SOS(846), BI=>SUB_BOS(877), OKI=>SUB_OKOS(879), BO=>SUB_BOS(878), OKO=>SUB_OKOS(878), D=>SUB_DS(878), SO=>SUB_SOS(878));
	DIV879: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(846), SI=>SUB_SOS(847), BI=>SUB_BOS(878), OKI=>SUB_OKOS(880), BO=>SUB_BOS(879), OKO=>SUB_OKOS(879), D=>SUB_DS(879), SO=>SUB_SOS(879));
	DIV880: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(847), SI=>SUB_SOS(848), BI=>SUB_BOS(879), OKI=>SUB_OKOS(881), BO=>SUB_BOS(880), OKO=>SUB_OKOS(880), D=>SUB_DS(880), SO=>SUB_SOS(880));
	DIV881: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(848), SI=>SUB_SOS(849), BI=>SUB_BOS(880), OKI=>SUB_OKOS(882), BO=>SUB_BOS(881), OKO=>SUB_OKOS(881), D=>SUB_DS(881), SO=>SUB_SOS(881));
	DIV882: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(849), SI=>SUB_SOS(850), BI=>SUB_BOS(881), OKI=>SUB_OKOS(883), BO=>SUB_BOS(882), OKO=>SUB_OKOS(882), D=>SUB_DS(882), SO=>SUB_SOS(882));
	DIV883: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(850), SI=>SUB_SOS(851), BI=>SUB_BOS(882), OKI=>SUB_OKOS(884), BO=>SUB_BOS(883), OKO=>SUB_OKOS(883), D=>SUB_DS(883), SO=>SUB_SOS(883));
	DIV884: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(851), SI=>SUB_SOS(852), BI=>SUB_BOS(883), OKI=>SUB_OKOS(885), BO=>SUB_BOS(884), OKO=>SUB_OKOS(884), D=>SUB_DS(884), SO=>SUB_SOS(884));
	DIV885: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(852), SI=>SUB_SOS(853), BI=>SUB_BOS(884), OKI=>SUB_OKOS(886), BO=>SUB_BOS(885), OKO=>SUB_OKOS(885), D=>SUB_DS(885), SO=>SUB_SOS(885));
	DIV886: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(853), SI=>SUB_SOS(854), BI=>SUB_BOS(885), OKI=>SUB_OKOS(887), BO=>SUB_BOS(886), OKO=>SUB_OKOS(886), D=>SUB_DS(886), SO=>SUB_SOS(886));
	DIV887: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(854), SI=>SUB_SOS(855), BI=>SUB_BOS(886), OKI=>SUB_OKOS(888), BO=>SUB_BOS(887), OKO=>SUB_OKOS(887), D=>SUB_DS(887), SO=>SUB_SOS(887));
	DIV888: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(855), SI=>SUB_SOS(856), BI=>SUB_BOS(887), OKI=>SUB_OKOS(889), BO=>SUB_BOS(888), OKO=>SUB_OKOS(888), D=>SUB_DS(888), SO=>SUB_SOS(888));
	DIV889: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(856), SI=>SUB_SOS(857), BI=>SUB_BOS(888), OKI=>SUB_OKOS(890), BO=>SUB_BOS(889), OKO=>SUB_OKOS(889), D=>SUB_DS(889), SO=>SUB_SOS(889));
	DIV890: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(857), SI=>SUB_SOS(858), BI=>SUB_BOS(889), OKI=>SUB_OKOS(891), BO=>SUB_BOS(890), OKO=>SUB_OKOS(890), D=>SUB_DS(890), SO=>SUB_SOS(890));
	DIV891: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(858), SI=>SUB_SOS(859), BI=>SUB_BOS(890), OKI=>SUB_OKOS(892), BO=>SUB_BOS(891), OKO=>SUB_OKOS(891), D=>SUB_DS(891), SO=>SUB_SOS(891));
	DIV892: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(859), SI=>SUB_SOS(860), BI=>SUB_BOS(891), OKI=>SUB_OKOS(893), BO=>SUB_BOS(892), OKO=>SUB_OKOS(892), D=>SUB_DS(892), SO=>SUB_SOS(892));
	DIV893: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(860), SI=>SUB_SOS(861), BI=>SUB_BOS(892), OKI=>SUB_OKOS(894), BO=>SUB_BOS(893), OKO=>SUB_OKOS(893), D=>SUB_DS(893), SO=>SUB_SOS(893));
	DIV894: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(861), SI=>SUB_SOS(862), BI=>SUB_BOS(893), OKI=>SUB_OKOS(895), BO=>SUB_BOS(894), OKO=>SUB_OKOS(894), D=>SUB_DS(894), SO=>SUB_SOS(894));
	DIV895: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(862), SI=>SUB_SOS(863), BI=>SUB_BOS(894), OKI=>BONS(27), BO=>SUB_BOS(895), OKO=>SUB_OKOS(895), D=>SUB_DS(895), SO=>SUB_SOS(895));

	DIV896: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(3), SI=>SUB_SOS(864), BI=>'0', OKI=>SUB_OKOS(897), BO=>SUB_BOS(896), OKO=>SUB_OKOS(896), D=>SUB_DS(896), SO=>SUB_SOS(896));
	DIV897: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(864), SI=>SUB_SOS(865), BI=>SUB_BOS(896), OKI=>SUB_OKOS(898), BO=>SUB_BOS(897), OKO=>SUB_OKOS(897), D=>SUB_DS(897), SO=>SUB_SOS(897));
	DIV898: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(865), SI=>SUB_SOS(866), BI=>SUB_BOS(897), OKI=>SUB_OKOS(899), BO=>SUB_BOS(898), OKO=>SUB_OKOS(898), D=>SUB_DS(898), SO=>SUB_SOS(898));
	DIV899: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(866), SI=>SUB_SOS(867), BI=>SUB_BOS(898), OKI=>SUB_OKOS(900), BO=>SUB_BOS(899), OKO=>SUB_OKOS(899), D=>SUB_DS(899), SO=>SUB_SOS(899));
	DIV900: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(867), SI=>SUB_SOS(868), BI=>SUB_BOS(899), OKI=>SUB_OKOS(901), BO=>SUB_BOS(900), OKO=>SUB_OKOS(900), D=>SUB_DS(900), SO=>SUB_SOS(900));
	DIV901: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(868), SI=>SUB_SOS(869), BI=>SUB_BOS(900), OKI=>SUB_OKOS(902), BO=>SUB_BOS(901), OKO=>SUB_OKOS(901), D=>SUB_DS(901), SO=>SUB_SOS(901));
	DIV902: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(869), SI=>SUB_SOS(870), BI=>SUB_BOS(901), OKI=>SUB_OKOS(903), BO=>SUB_BOS(902), OKO=>SUB_OKOS(902), D=>SUB_DS(902), SO=>SUB_SOS(902));
	DIV903: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(870), SI=>SUB_SOS(871), BI=>SUB_BOS(902), OKI=>SUB_OKOS(904), BO=>SUB_BOS(903), OKO=>SUB_OKOS(903), D=>SUB_DS(903), SO=>SUB_SOS(903));
	DIV904: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(871), SI=>SUB_SOS(872), BI=>SUB_BOS(903), OKI=>SUB_OKOS(905), BO=>SUB_BOS(904), OKO=>SUB_OKOS(904), D=>SUB_DS(904), SO=>SUB_SOS(904));
	DIV905: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(872), SI=>SUB_SOS(873), BI=>SUB_BOS(904), OKI=>SUB_OKOS(906), BO=>SUB_BOS(905), OKO=>SUB_OKOS(905), D=>SUB_DS(905), SO=>SUB_SOS(905));
	DIV906: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(873), SI=>SUB_SOS(874), BI=>SUB_BOS(905), OKI=>SUB_OKOS(907), BO=>SUB_BOS(906), OKO=>SUB_OKOS(906), D=>SUB_DS(906), SO=>SUB_SOS(906));
	DIV907: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(874), SI=>SUB_SOS(875), BI=>SUB_BOS(906), OKI=>SUB_OKOS(908), BO=>SUB_BOS(907), OKO=>SUB_OKOS(907), D=>SUB_DS(907), SO=>SUB_SOS(907));
	DIV908: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(875), SI=>SUB_SOS(876), BI=>SUB_BOS(907), OKI=>SUB_OKOS(909), BO=>SUB_BOS(908), OKO=>SUB_OKOS(908), D=>SUB_DS(908), SO=>SUB_SOS(908));
	DIV909: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(876), SI=>SUB_SOS(877), BI=>SUB_BOS(908), OKI=>SUB_OKOS(910), BO=>SUB_BOS(909), OKO=>SUB_OKOS(909), D=>SUB_DS(909), SO=>SUB_SOS(909));
	DIV910: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(877), SI=>SUB_SOS(878), BI=>SUB_BOS(909), OKI=>SUB_OKOS(911), BO=>SUB_BOS(910), OKO=>SUB_OKOS(910), D=>SUB_DS(910), SO=>SUB_SOS(910));
	DIV911: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(878), SI=>SUB_SOS(879), BI=>SUB_BOS(910), OKI=>SUB_OKOS(912), BO=>SUB_BOS(911), OKO=>SUB_OKOS(911), D=>SUB_DS(911), SO=>SUB_SOS(911));
	DIV912: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(879), SI=>SUB_SOS(880), BI=>SUB_BOS(911), OKI=>SUB_OKOS(913), BO=>SUB_BOS(912), OKO=>SUB_OKOS(912), D=>SUB_DS(912), SO=>SUB_SOS(912));
	DIV913: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(880), SI=>SUB_SOS(881), BI=>SUB_BOS(912), OKI=>SUB_OKOS(914), BO=>SUB_BOS(913), OKO=>SUB_OKOS(913), D=>SUB_DS(913), SO=>SUB_SOS(913));
	DIV914: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(881), SI=>SUB_SOS(882), BI=>SUB_BOS(913), OKI=>SUB_OKOS(915), BO=>SUB_BOS(914), OKO=>SUB_OKOS(914), D=>SUB_DS(914), SO=>SUB_SOS(914));
	DIV915: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(882), SI=>SUB_SOS(883), BI=>SUB_BOS(914), OKI=>SUB_OKOS(916), BO=>SUB_BOS(915), OKO=>SUB_OKOS(915), D=>SUB_DS(915), SO=>SUB_SOS(915));
	DIV916: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(883), SI=>SUB_SOS(884), BI=>SUB_BOS(915), OKI=>SUB_OKOS(917), BO=>SUB_BOS(916), OKO=>SUB_OKOS(916), D=>SUB_DS(916), SO=>SUB_SOS(916));
	DIV917: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(884), SI=>SUB_SOS(885), BI=>SUB_BOS(916), OKI=>SUB_OKOS(918), BO=>SUB_BOS(917), OKO=>SUB_OKOS(917), D=>SUB_DS(917), SO=>SUB_SOS(917));
	DIV918: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(885), SI=>SUB_SOS(886), BI=>SUB_BOS(917), OKI=>SUB_OKOS(919), BO=>SUB_BOS(918), OKO=>SUB_OKOS(918), D=>SUB_DS(918), SO=>SUB_SOS(918));
	DIV919: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(886), SI=>SUB_SOS(887), BI=>SUB_BOS(918), OKI=>SUB_OKOS(920), BO=>SUB_BOS(919), OKO=>SUB_OKOS(919), D=>SUB_DS(919), SO=>SUB_SOS(919));
	DIV920: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(887), SI=>SUB_SOS(888), BI=>SUB_BOS(919), OKI=>SUB_OKOS(921), BO=>SUB_BOS(920), OKO=>SUB_OKOS(920), D=>SUB_DS(920), SO=>SUB_SOS(920));
	DIV921: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(888), SI=>SUB_SOS(889), BI=>SUB_BOS(920), OKI=>SUB_OKOS(922), BO=>SUB_BOS(921), OKO=>SUB_OKOS(921), D=>SUB_DS(921), SO=>SUB_SOS(921));
	DIV922: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(889), SI=>SUB_SOS(890), BI=>SUB_BOS(921), OKI=>SUB_OKOS(923), BO=>SUB_BOS(922), OKO=>SUB_OKOS(922), D=>SUB_DS(922), SO=>SUB_SOS(922));
	DIV923: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(890), SI=>SUB_SOS(891), BI=>SUB_BOS(922), OKI=>SUB_OKOS(924), BO=>SUB_BOS(923), OKO=>SUB_OKOS(923), D=>SUB_DS(923), SO=>SUB_SOS(923));
	DIV924: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(891), SI=>SUB_SOS(892), BI=>SUB_BOS(923), OKI=>SUB_OKOS(925), BO=>SUB_BOS(924), OKO=>SUB_OKOS(924), D=>SUB_DS(924), SO=>SUB_SOS(924));
	DIV925: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(892), SI=>SUB_SOS(893), BI=>SUB_BOS(924), OKI=>SUB_OKOS(926), BO=>SUB_BOS(925), OKO=>SUB_OKOS(925), D=>SUB_DS(925), SO=>SUB_SOS(925));
	DIV926: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(893), SI=>SUB_SOS(894), BI=>SUB_BOS(925), OKI=>SUB_OKOS(927), BO=>SUB_BOS(926), OKO=>SUB_OKOS(926), D=>SUB_DS(926), SO=>SUB_SOS(926));
	DIV927: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(894), SI=>SUB_SOS(895), BI=>SUB_BOS(926), OKI=>BONS(28), BO=>SUB_BOS(927), OKO=>SUB_OKOS(927), D=>SUB_DS(927), SO=>SUB_SOS(927));

	DIV928: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(2), SI=>SUB_SOS(896), BI=>'0', OKI=>SUB_OKOS(929), BO=>SUB_BOS(928), OKO=>SUB_OKOS(928), D=>SUB_DS(928), SO=>SUB_SOS(928));
	DIV929: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(896), SI=>SUB_SOS(897), BI=>SUB_BOS(928), OKI=>SUB_OKOS(930), BO=>SUB_BOS(929), OKO=>SUB_OKOS(929), D=>SUB_DS(929), SO=>SUB_SOS(929));
	DIV930: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(897), SI=>SUB_SOS(898), BI=>SUB_BOS(929), OKI=>SUB_OKOS(931), BO=>SUB_BOS(930), OKO=>SUB_OKOS(930), D=>SUB_DS(930), SO=>SUB_SOS(930));
	DIV931: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(898), SI=>SUB_SOS(899), BI=>SUB_BOS(930), OKI=>SUB_OKOS(932), BO=>SUB_BOS(931), OKO=>SUB_OKOS(931), D=>SUB_DS(931), SO=>SUB_SOS(931));
	DIV932: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(899), SI=>SUB_SOS(900), BI=>SUB_BOS(931), OKI=>SUB_OKOS(933), BO=>SUB_BOS(932), OKO=>SUB_OKOS(932), D=>SUB_DS(932), SO=>SUB_SOS(932));
	DIV933: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(900), SI=>SUB_SOS(901), BI=>SUB_BOS(932), OKI=>SUB_OKOS(934), BO=>SUB_BOS(933), OKO=>SUB_OKOS(933), D=>SUB_DS(933), SO=>SUB_SOS(933));
	DIV934: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(901), SI=>SUB_SOS(902), BI=>SUB_BOS(933), OKI=>SUB_OKOS(935), BO=>SUB_BOS(934), OKO=>SUB_OKOS(934), D=>SUB_DS(934), SO=>SUB_SOS(934));
	DIV935: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(902), SI=>SUB_SOS(903), BI=>SUB_BOS(934), OKI=>SUB_OKOS(936), BO=>SUB_BOS(935), OKO=>SUB_OKOS(935), D=>SUB_DS(935), SO=>SUB_SOS(935));
	DIV936: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(903), SI=>SUB_SOS(904), BI=>SUB_BOS(935), OKI=>SUB_OKOS(937), BO=>SUB_BOS(936), OKO=>SUB_OKOS(936), D=>SUB_DS(936), SO=>SUB_SOS(936));
	DIV937: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(904), SI=>SUB_SOS(905), BI=>SUB_BOS(936), OKI=>SUB_OKOS(938), BO=>SUB_BOS(937), OKO=>SUB_OKOS(937), D=>SUB_DS(937), SO=>SUB_SOS(937));
	DIV938: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(905), SI=>SUB_SOS(906), BI=>SUB_BOS(937), OKI=>SUB_OKOS(939), BO=>SUB_BOS(938), OKO=>SUB_OKOS(938), D=>SUB_DS(938), SO=>SUB_SOS(938));
	DIV939: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(906), SI=>SUB_SOS(907), BI=>SUB_BOS(938), OKI=>SUB_OKOS(940), BO=>SUB_BOS(939), OKO=>SUB_OKOS(939), D=>SUB_DS(939), SO=>SUB_SOS(939));
	DIV940: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(907), SI=>SUB_SOS(908), BI=>SUB_BOS(939), OKI=>SUB_OKOS(941), BO=>SUB_BOS(940), OKO=>SUB_OKOS(940), D=>SUB_DS(940), SO=>SUB_SOS(940));
	DIV941: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(908), SI=>SUB_SOS(909), BI=>SUB_BOS(940), OKI=>SUB_OKOS(942), BO=>SUB_BOS(941), OKO=>SUB_OKOS(941), D=>SUB_DS(941), SO=>SUB_SOS(941));
	DIV942: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(909), SI=>SUB_SOS(910), BI=>SUB_BOS(941), OKI=>SUB_OKOS(943), BO=>SUB_BOS(942), OKO=>SUB_OKOS(942), D=>SUB_DS(942), SO=>SUB_SOS(942));
	DIV943: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(910), SI=>SUB_SOS(911), BI=>SUB_BOS(942), OKI=>SUB_OKOS(944), BO=>SUB_BOS(943), OKO=>SUB_OKOS(943), D=>SUB_DS(943), SO=>SUB_SOS(943));
	DIV944: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(911), SI=>SUB_SOS(912), BI=>SUB_BOS(943), OKI=>SUB_OKOS(945), BO=>SUB_BOS(944), OKO=>SUB_OKOS(944), D=>SUB_DS(944), SO=>SUB_SOS(944));
	DIV945: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(912), SI=>SUB_SOS(913), BI=>SUB_BOS(944), OKI=>SUB_OKOS(946), BO=>SUB_BOS(945), OKO=>SUB_OKOS(945), D=>SUB_DS(945), SO=>SUB_SOS(945));
	DIV946: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(913), SI=>SUB_SOS(914), BI=>SUB_BOS(945), OKI=>SUB_OKOS(947), BO=>SUB_BOS(946), OKO=>SUB_OKOS(946), D=>SUB_DS(946), SO=>SUB_SOS(946));
	DIV947: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(914), SI=>SUB_SOS(915), BI=>SUB_BOS(946), OKI=>SUB_OKOS(948), BO=>SUB_BOS(947), OKO=>SUB_OKOS(947), D=>SUB_DS(947), SO=>SUB_SOS(947));
	DIV948: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(915), SI=>SUB_SOS(916), BI=>SUB_BOS(947), OKI=>SUB_OKOS(949), BO=>SUB_BOS(948), OKO=>SUB_OKOS(948), D=>SUB_DS(948), SO=>SUB_SOS(948));
	DIV949: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(916), SI=>SUB_SOS(917), BI=>SUB_BOS(948), OKI=>SUB_OKOS(950), BO=>SUB_BOS(949), OKO=>SUB_OKOS(949), D=>SUB_DS(949), SO=>SUB_SOS(949));
	DIV950: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(917), SI=>SUB_SOS(918), BI=>SUB_BOS(949), OKI=>SUB_OKOS(951), BO=>SUB_BOS(950), OKO=>SUB_OKOS(950), D=>SUB_DS(950), SO=>SUB_SOS(950));
	DIV951: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(918), SI=>SUB_SOS(919), BI=>SUB_BOS(950), OKI=>SUB_OKOS(952), BO=>SUB_BOS(951), OKO=>SUB_OKOS(951), D=>SUB_DS(951), SO=>SUB_SOS(951));
	DIV952: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(919), SI=>SUB_SOS(920), BI=>SUB_BOS(951), OKI=>SUB_OKOS(953), BO=>SUB_BOS(952), OKO=>SUB_OKOS(952), D=>SUB_DS(952), SO=>SUB_SOS(952));
	DIV953: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(920), SI=>SUB_SOS(921), BI=>SUB_BOS(952), OKI=>SUB_OKOS(954), BO=>SUB_BOS(953), OKO=>SUB_OKOS(953), D=>SUB_DS(953), SO=>SUB_SOS(953));
	DIV954: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(921), SI=>SUB_SOS(922), BI=>SUB_BOS(953), OKI=>SUB_OKOS(955), BO=>SUB_BOS(954), OKO=>SUB_OKOS(954), D=>SUB_DS(954), SO=>SUB_SOS(954));
	DIV955: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(922), SI=>SUB_SOS(923), BI=>SUB_BOS(954), OKI=>SUB_OKOS(956), BO=>SUB_BOS(955), OKO=>SUB_OKOS(955), D=>SUB_DS(955), SO=>SUB_SOS(955));
	DIV956: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(923), SI=>SUB_SOS(924), BI=>SUB_BOS(955), OKI=>SUB_OKOS(957), BO=>SUB_BOS(956), OKO=>SUB_OKOS(956), D=>SUB_DS(956), SO=>SUB_SOS(956));
	DIV957: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(924), SI=>SUB_SOS(925), BI=>SUB_BOS(956), OKI=>SUB_OKOS(958), BO=>SUB_BOS(957), OKO=>SUB_OKOS(957), D=>SUB_DS(957), SO=>SUB_SOS(957));
	DIV958: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(925), SI=>SUB_SOS(926), BI=>SUB_BOS(957), OKI=>SUB_OKOS(959), BO=>SUB_BOS(958), OKO=>SUB_OKOS(958), D=>SUB_DS(958), SO=>SUB_SOS(958));
	DIV959: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(926), SI=>SUB_SOS(927), BI=>SUB_BOS(958), OKI=>BONS(29), BO=>SUB_BOS(959), OKO=>SUB_OKOS(959), D=>SUB_DS(959), SO=>SUB_SOS(959));

	DIV960: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(1), SI=>SUB_SOS(928), BI=>'0', OKI=>SUB_OKOS(961), BO=>SUB_BOS(960), OKO=>SUB_OKOS(960), D=>SUB_DS(960), SO=>SUB_SOS(960));
	DIV961: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(928), SI=>SUB_SOS(929), BI=>SUB_BOS(960), OKI=>SUB_OKOS(962), BO=>SUB_BOS(961), OKO=>SUB_OKOS(961), D=>SUB_DS(961), SO=>SUB_SOS(961));
	DIV962: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(929), SI=>SUB_SOS(930), BI=>SUB_BOS(961), OKI=>SUB_OKOS(963), BO=>SUB_BOS(962), OKO=>SUB_OKOS(962), D=>SUB_DS(962), SO=>SUB_SOS(962));
	DIV963: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(930), SI=>SUB_SOS(931), BI=>SUB_BOS(962), OKI=>SUB_OKOS(964), BO=>SUB_BOS(963), OKO=>SUB_OKOS(963), D=>SUB_DS(963), SO=>SUB_SOS(963));
	DIV964: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(931), SI=>SUB_SOS(932), BI=>SUB_BOS(963), OKI=>SUB_OKOS(965), BO=>SUB_BOS(964), OKO=>SUB_OKOS(964), D=>SUB_DS(964), SO=>SUB_SOS(964));
	DIV965: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(932), SI=>SUB_SOS(933), BI=>SUB_BOS(964), OKI=>SUB_OKOS(966), BO=>SUB_BOS(965), OKO=>SUB_OKOS(965), D=>SUB_DS(965), SO=>SUB_SOS(965));
	DIV966: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(933), SI=>SUB_SOS(934), BI=>SUB_BOS(965), OKI=>SUB_OKOS(967), BO=>SUB_BOS(966), OKO=>SUB_OKOS(966), D=>SUB_DS(966), SO=>SUB_SOS(966));
	DIV967: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(934), SI=>SUB_SOS(935), BI=>SUB_BOS(966), OKI=>SUB_OKOS(968), BO=>SUB_BOS(967), OKO=>SUB_OKOS(967), D=>SUB_DS(967), SO=>SUB_SOS(967));
	DIV968: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(935), SI=>SUB_SOS(936), BI=>SUB_BOS(967), OKI=>SUB_OKOS(969), BO=>SUB_BOS(968), OKO=>SUB_OKOS(968), D=>SUB_DS(968), SO=>SUB_SOS(968));
	DIV969: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(936), SI=>SUB_SOS(937), BI=>SUB_BOS(968), OKI=>SUB_OKOS(970), BO=>SUB_BOS(969), OKO=>SUB_OKOS(969), D=>SUB_DS(969), SO=>SUB_SOS(969));
	DIV970: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(937), SI=>SUB_SOS(938), BI=>SUB_BOS(969), OKI=>SUB_OKOS(971), BO=>SUB_BOS(970), OKO=>SUB_OKOS(970), D=>SUB_DS(970), SO=>SUB_SOS(970));
	DIV971: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(938), SI=>SUB_SOS(939), BI=>SUB_BOS(970), OKI=>SUB_OKOS(972), BO=>SUB_BOS(971), OKO=>SUB_OKOS(971), D=>SUB_DS(971), SO=>SUB_SOS(971));
	DIV972: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(939), SI=>SUB_SOS(940), BI=>SUB_BOS(971), OKI=>SUB_OKOS(973), BO=>SUB_BOS(972), OKO=>SUB_OKOS(972), D=>SUB_DS(972), SO=>SUB_SOS(972));
	DIV973: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(940), SI=>SUB_SOS(941), BI=>SUB_BOS(972), OKI=>SUB_OKOS(974), BO=>SUB_BOS(973), OKO=>SUB_OKOS(973), D=>SUB_DS(973), SO=>SUB_SOS(973));
	DIV974: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(941), SI=>SUB_SOS(942), BI=>SUB_BOS(973), OKI=>SUB_OKOS(975), BO=>SUB_BOS(974), OKO=>SUB_OKOS(974), D=>SUB_DS(974), SO=>SUB_SOS(974));
	DIV975: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(942), SI=>SUB_SOS(943), BI=>SUB_BOS(974), OKI=>SUB_OKOS(976), BO=>SUB_BOS(975), OKO=>SUB_OKOS(975), D=>SUB_DS(975), SO=>SUB_SOS(975));
	DIV976: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(943), SI=>SUB_SOS(944), BI=>SUB_BOS(975), OKI=>SUB_OKOS(977), BO=>SUB_BOS(976), OKO=>SUB_OKOS(976), D=>SUB_DS(976), SO=>SUB_SOS(976));
	DIV977: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(944), SI=>SUB_SOS(945), BI=>SUB_BOS(976), OKI=>SUB_OKOS(978), BO=>SUB_BOS(977), OKO=>SUB_OKOS(977), D=>SUB_DS(977), SO=>SUB_SOS(977));
	DIV978: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(945), SI=>SUB_SOS(946), BI=>SUB_BOS(977), OKI=>SUB_OKOS(979), BO=>SUB_BOS(978), OKO=>SUB_OKOS(978), D=>SUB_DS(978), SO=>SUB_SOS(978));
	DIV979: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(946), SI=>SUB_SOS(947), BI=>SUB_BOS(978), OKI=>SUB_OKOS(980), BO=>SUB_BOS(979), OKO=>SUB_OKOS(979), D=>SUB_DS(979), SO=>SUB_SOS(979));
	DIV980: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(947), SI=>SUB_SOS(948), BI=>SUB_BOS(979), OKI=>SUB_OKOS(981), BO=>SUB_BOS(980), OKO=>SUB_OKOS(980), D=>SUB_DS(980), SO=>SUB_SOS(980));
	DIV981: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(948), SI=>SUB_SOS(949), BI=>SUB_BOS(980), OKI=>SUB_OKOS(982), BO=>SUB_BOS(981), OKO=>SUB_OKOS(981), D=>SUB_DS(981), SO=>SUB_SOS(981));
	DIV982: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(949), SI=>SUB_SOS(950), BI=>SUB_BOS(981), OKI=>SUB_OKOS(983), BO=>SUB_BOS(982), OKO=>SUB_OKOS(982), D=>SUB_DS(982), SO=>SUB_SOS(982));
	DIV983: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(950), SI=>SUB_SOS(951), BI=>SUB_BOS(982), OKI=>SUB_OKOS(984), BO=>SUB_BOS(983), OKO=>SUB_OKOS(983), D=>SUB_DS(983), SO=>SUB_SOS(983));
	DIV984: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(951), SI=>SUB_SOS(952), BI=>SUB_BOS(983), OKI=>SUB_OKOS(985), BO=>SUB_BOS(984), OKO=>SUB_OKOS(984), D=>SUB_DS(984), SO=>SUB_SOS(984));
	DIV985: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(952), SI=>SUB_SOS(953), BI=>SUB_BOS(984), OKI=>SUB_OKOS(986), BO=>SUB_BOS(985), OKO=>SUB_OKOS(985), D=>SUB_DS(985), SO=>SUB_SOS(985));
	DIV986: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(953), SI=>SUB_SOS(954), BI=>SUB_BOS(985), OKI=>SUB_OKOS(987), BO=>SUB_BOS(986), OKO=>SUB_OKOS(986), D=>SUB_DS(986), SO=>SUB_SOS(986));
	DIV987: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(954), SI=>SUB_SOS(955), BI=>SUB_BOS(986), OKI=>SUB_OKOS(988), BO=>SUB_BOS(987), OKO=>SUB_OKOS(987), D=>SUB_DS(987), SO=>SUB_SOS(987));
	DIV988: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(955), SI=>SUB_SOS(956), BI=>SUB_BOS(987), OKI=>SUB_OKOS(989), BO=>SUB_BOS(988), OKO=>SUB_OKOS(988), D=>SUB_DS(988), SO=>SUB_SOS(988));
	DIV989: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(956), SI=>SUB_SOS(957), BI=>SUB_BOS(988), OKI=>SUB_OKOS(990), BO=>SUB_BOS(989), OKO=>SUB_OKOS(989), D=>SUB_DS(989), SO=>SUB_SOS(989));
	DIV990: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(957), SI=>SUB_SOS(958), BI=>SUB_BOS(989), OKI=>SUB_OKOS(991), BO=>SUB_BOS(990), OKO=>SUB_OKOS(990), D=>SUB_DS(990), SO=>SUB_SOS(990));
	DIV991: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(958), SI=>SUB_SOS(959), BI=>SUB_BOS(990), OKI=>BONS(30), BO=>SUB_BOS(991), OKO=>SUB_OKOS(991), D=>SUB_DS(991), SO=>SUB_SOS(991));

	DIV992: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>DIVIDEND(0), SI=>SUB_SOS(960), BI=>'0', OKI=>SUB_OKOS(993), BO=>SUB_BOS(992), OKO=>SUB_OKOS(992), D=>SUB_DS(992), SO=>SUB_SOS(992));
	DIV993: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(960), SI=>SUB_SOS(961), BI=>SUB_BOS(992), OKI=>SUB_OKOS(994), BO=>SUB_BOS(993), OKO=>SUB_OKOS(993), D=>SUB_DS(993), SO=>SUB_SOS(993));
	DIV994: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(961), SI=>SUB_SOS(962), BI=>SUB_BOS(993), OKI=>SUB_OKOS(995), BO=>SUB_BOS(994), OKO=>SUB_OKOS(994), D=>SUB_DS(994), SO=>SUB_SOS(994));
	DIV995: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(962), SI=>SUB_SOS(963), BI=>SUB_BOS(994), OKI=>SUB_OKOS(996), BO=>SUB_BOS(995), OKO=>SUB_OKOS(995), D=>SUB_DS(995), SO=>SUB_SOS(995));
	DIV996: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(963), SI=>SUB_SOS(964), BI=>SUB_BOS(995), OKI=>SUB_OKOS(997), BO=>SUB_BOS(996), OKO=>SUB_OKOS(996), D=>SUB_DS(996), SO=>SUB_SOS(996));
	DIV997: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(964), SI=>SUB_SOS(965), BI=>SUB_BOS(996), OKI=>SUB_OKOS(998), BO=>SUB_BOS(997), OKO=>SUB_OKOS(997), D=>SUB_DS(997), SO=>SUB_SOS(997));
	DIV998: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(965), SI=>SUB_SOS(966), BI=>SUB_BOS(997), OKI=>SUB_OKOS(999), BO=>SUB_BOS(998), OKO=>SUB_OKOS(998), D=>SUB_DS(998), SO=>SUB_SOS(998));
	DIV999: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(966), SI=>SUB_SOS(967), BI=>SUB_BOS(998), OKI=>SUB_OKOS(1000), BO=>SUB_BOS(999), OKO=>SUB_OKOS(999), D=>SUB_DS(999), SO=>SUB_SOS(999));
	DIV1000: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(967), SI=>SUB_SOS(968), BI=>SUB_BOS(999), OKI=>SUB_OKOS(1001), BO=>SUB_BOS(1000), OKO=>SUB_OKOS(1000), D=>SUB_DS(1000), SO=>SUB_SOS(1000));
	DIV1001: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(968), SI=>SUB_SOS(969), BI=>SUB_BOS(1000), OKI=>SUB_OKOS(1002), BO=>SUB_BOS(1001), OKO=>SUB_OKOS(1001), D=>SUB_DS(1001), SO=>SUB_SOS(1001));
	DIV1002: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(969), SI=>SUB_SOS(970), BI=>SUB_BOS(1001), OKI=>SUB_OKOS(1003), BO=>SUB_BOS(1002), OKO=>SUB_OKOS(1002), D=>SUB_DS(1002), SO=>SUB_SOS(1002));
	DIV1003: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(970), SI=>SUB_SOS(971), BI=>SUB_BOS(1002), OKI=>SUB_OKOS(1004), BO=>SUB_BOS(1003), OKO=>SUB_OKOS(1003), D=>SUB_DS(1003), SO=>SUB_SOS(1003));
	DIV1004: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(971), SI=>SUB_SOS(972), BI=>SUB_BOS(1003), OKI=>SUB_OKOS(1005), BO=>SUB_BOS(1004), OKO=>SUB_OKOS(1004), D=>SUB_DS(1004), SO=>SUB_SOS(1004));
	DIV1005: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(972), SI=>SUB_SOS(973), BI=>SUB_BOS(1004), OKI=>SUB_OKOS(1006), BO=>SUB_BOS(1005), OKO=>SUB_OKOS(1005), D=>SUB_DS(1005), SO=>SUB_SOS(1005));
	DIV1006: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(973), SI=>SUB_SOS(974), BI=>SUB_BOS(1005), OKI=>SUB_OKOS(1007), BO=>SUB_BOS(1006), OKO=>SUB_OKOS(1006), D=>SUB_DS(1006), SO=>SUB_SOS(1006));
	DIV1007: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(974), SI=>SUB_SOS(975), BI=>SUB_BOS(1006), OKI=>SUB_OKOS(1008), BO=>SUB_BOS(1007), OKO=>SUB_OKOS(1007), D=>SUB_DS(1007), SO=>SUB_SOS(1007));
	DIV1008: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(975), SI=>SUB_SOS(976), BI=>SUB_BOS(1007), OKI=>SUB_OKOS(1009), BO=>SUB_BOS(1008), OKO=>SUB_OKOS(1008), D=>SUB_DS(1008), SO=>SUB_SOS(1008));
	DIV1009: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(976), SI=>SUB_SOS(977), BI=>SUB_BOS(1008), OKI=>SUB_OKOS(1010), BO=>SUB_BOS(1009), OKO=>SUB_OKOS(1009), D=>SUB_DS(1009), SO=>SUB_SOS(1009));
	DIV1010: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(977), SI=>SUB_SOS(978), BI=>SUB_BOS(1009), OKI=>SUB_OKOS(1011), BO=>SUB_BOS(1010), OKO=>SUB_OKOS(1010), D=>SUB_DS(1010), SO=>SUB_SOS(1010));
	DIV1011: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(978), SI=>SUB_SOS(979), BI=>SUB_BOS(1010), OKI=>SUB_OKOS(1012), BO=>SUB_BOS(1011), OKO=>SUB_OKOS(1011), D=>SUB_DS(1011), SO=>SUB_SOS(1011));
	DIV1012: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(979), SI=>SUB_SOS(980), BI=>SUB_BOS(1011), OKI=>SUB_OKOS(1013), BO=>SUB_BOS(1012), OKO=>SUB_OKOS(1012), D=>SUB_DS(1012), SO=>SUB_SOS(1012));
	DIV1013: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(980), SI=>SUB_SOS(981), BI=>SUB_BOS(1012), OKI=>SUB_OKOS(1014), BO=>SUB_BOS(1013), OKO=>SUB_OKOS(1013), D=>SUB_DS(1013), SO=>SUB_SOS(1013));
	DIV1014: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(981), SI=>SUB_SOS(982), BI=>SUB_BOS(1013), OKI=>SUB_OKOS(1015), BO=>SUB_BOS(1014), OKO=>SUB_OKOS(1014), D=>SUB_DS(1014), SO=>SUB_SOS(1014));
	DIV1015: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(982), SI=>SUB_SOS(983), BI=>SUB_BOS(1014), OKI=>SUB_OKOS(1016), BO=>SUB_BOS(1015), OKO=>SUB_OKOS(1015), D=>SUB_DS(1015), SO=>SUB_SOS(1015));
	DIV1016: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(983), SI=>SUB_SOS(984), BI=>SUB_BOS(1015), OKI=>SUB_OKOS(1017), BO=>SUB_BOS(1016), OKO=>SUB_OKOS(1016), D=>SUB_DS(1016), SO=>SUB_SOS(1016));
	DIV1017: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(984), SI=>SUB_SOS(985), BI=>SUB_BOS(1016), OKI=>SUB_OKOS(1018), BO=>SUB_BOS(1017), OKO=>SUB_OKOS(1017), D=>SUB_DS(1017), SO=>SUB_SOS(1017));
	DIV1018: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(985), SI=>SUB_SOS(986), BI=>SUB_BOS(1017), OKI=>SUB_OKOS(1019), BO=>SUB_BOS(1018), OKO=>SUB_OKOS(1018), D=>SUB_DS(1018), SO=>SUB_SOS(1018));
	DIV1019: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(986), SI=>SUB_SOS(987), BI=>SUB_BOS(1018), OKI=>SUB_OKOS(1020), BO=>SUB_BOS(1019), OKO=>SUB_OKOS(1019), D=>SUB_DS(1019), SO=>SUB_SOS(1019));
	DIV1020: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(987), SI=>SUB_SOS(988), BI=>SUB_BOS(1019), OKI=>SUB_OKOS(1021), BO=>SUB_BOS(1020), OKO=>SUB_OKOS(1020), D=>SUB_DS(1020), SO=>SUB_SOS(1020));
	DIV1021: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(988), SI=>SUB_SOS(989), BI=>SUB_BOS(1020), OKI=>SUB_OKOS(1022), BO=>SUB_BOS(1021), OKO=>SUB_OKOS(1021), D=>SUB_DS(1021), SO=>SUB_SOS(1021));
	DIV1022: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(989), SI=>SUB_SOS(990), BI=>SUB_BOS(1021), OKI=>SUB_OKOS(1023), BO=>SUB_BOS(1022), OKO=>SUB_OKOS(1022), D=>SUB_DS(1022), SO=>SUB_SOS(1022));
	DIV1023: Chowdhury_1BitDiv_Dec7 PORT MAP(M=>SUB_DS(990), SI=>SUB_SOS(991), BI=>SUB_BOS(1022), OKI=>BONS(31), BO=>SUB_BOS(1023), OKO=>SUB_OKOS(1023), D=>SUB_DS(1023), SO=>SUB_SOS(1023));

	Q(0) <= SUB_OKOS(992);
	Q(1) <= SUB_OKOS(960);
	Q(2) <= SUB_OKOS(928);
	Q(3) <= SUB_OKOS(896);
	Q(4) <= SUB_OKOS(864);
	Q(5) <= SUB_OKOS(832);
	Q(6) <= SUB_OKOS(800);
	Q(7) <= SUB_OKOS(768);
	Q(8) <= SUB_OKOS(736);
	Q(9) <= SUB_OKOS(704);
	Q(10) <= SUB_OKOS(672);
	Q(11) <= SUB_OKOS(640);
	Q(12) <= SUB_OKOS(608);
	Q(13) <= SUB_OKOS(576);
	Q(14) <= SUB_OKOS(544);
	Q(15) <= SUB_OKOS(512);
	Q(16) <= SUB_OKOS(480);
	Q(17) <= SUB_OKOS(448);
	Q(18) <= SUB_OKOS(416);
	Q(19) <= SUB_OKOS(384);
	Q(20) <= SUB_OKOS(352);
	Q(21) <= SUB_OKOS(320);
	Q(22) <= SUB_OKOS(288);
	Q(23) <= SUB_OKOS(256);
	Q(24) <= SUB_OKOS(224);
	Q(25) <= SUB_OKOS(192);
	Q(26) <= SUB_OKOS(160);
	Q(27) <= SUB_OKOS(128);
	Q(28) <= SUB_OKOS(96);
	Q(29) <= SUB_OKOS(64);
	Q(30) <= SUB_OKOS(32);
	Q(31) <= SUB_OKOS(0);

	R(0) <= SUB_DS(992);
	R(1) <= SUB_DS(993);
	R(2) <= SUB_DS(994);
	R(3) <= SUB_DS(995);
	R(4) <= SUB_DS(996);
	R(5) <= SUB_DS(997);
	R(6) <= SUB_DS(998);
	R(7) <= SUB_DS(999);
	R(8) <= SUB_DS(1000);
	R(9) <= SUB_DS(1001);
	R(10) <= SUB_DS(1002);
	R(11) <= SUB_DS(1003);
	R(12) <= SUB_DS(1004);
	R(13) <= SUB_DS(1005);
	R(14) <= SUB_DS(1006);
	R(15) <= SUB_DS(1007);
	R(16) <= SUB_DS(1008);
	R(17) <= SUB_DS(1009);
	R(18) <= SUB_DS(1010);
	R(19) <= SUB_DS(1011);
	R(20) <= SUB_DS(1012);
	R(21) <= SUB_DS(1013);
	R(22) <= SUB_DS(1014);
	R(23) <= SUB_DS(1015);
	R(24) <= SUB_DS(1016);
	R(25) <= SUB_DS(1017);
	R(26) <= SUB_DS(1018);
	R(27) <= SUB_DS(1019);
	R(28) <= SUB_DS(1020);
	R(29) <= SUB_DS(1021);
	R(30) <= SUB_DS(1022);
	R(31) <= SUB_DS(1023);
	
	
	QUOTIENT <= Q;
	REMAINDER <= R;
	
END Chowdhury_Behaviour;