-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_MUX 

-- ============================================================
-- File Name: Chowdhury_LPM_32Bit64x1Mux_Dec7.vhd
-- Megafunction Name(s):
-- 			LPM_MUX
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 16.0.0 Build 211 04/27/2016 SJ Lite Edition
-- ************************************************************


--Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus Prime License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY Chowdhury_LPM_32Bit64x1Mux_Dec7 IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data10x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data11x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data12x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data13x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data14x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data15x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data16x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data17x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data18x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data19x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data20x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data21x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data22x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data23x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data24x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data25x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data26x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data27x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data28x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data29x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data30x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data31x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data32x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data33x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data34x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data35x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data36x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data37x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data38x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data39x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data40x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data41x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data42x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data43x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data44x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data45x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data46x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data47x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data48x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data49x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data50x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data51x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data52x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data53x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data54x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data55x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data56x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data57x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data58x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data59x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data60x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data61x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data62x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data63x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data8x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data9x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END Chowdhury_LPM_32Bit64x1Mux_Dec7;


ARCHITECTURE SYN OF chowdhury_lpm_32bit64x1mux_dec7 IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_2D (63 DOWNTO 0, 31 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire18	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire19	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire20	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire21	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire22	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire23	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire24	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire25	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire26	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire27	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire28	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire29	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire30	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire31	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire32	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire33	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire34	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire35	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire36	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire37	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire38	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire39	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire40	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire41	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire42	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire43	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire44	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire45	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire46	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire47	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire48	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire49	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire50	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire51	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire52	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire53	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire54	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire55	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire56	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire57	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire58	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire59	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire60	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire61	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire62	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire63	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire64	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire65	: STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
	sub_wire64    <= data0x(31 DOWNTO 0);
	sub_wire63    <= data1x(31 DOWNTO 0);
	sub_wire62    <= data2x(31 DOWNTO 0);
	sub_wire61    <= data3x(31 DOWNTO 0);
	sub_wire60    <= data4x(31 DOWNTO 0);
	sub_wire59    <= data5x(31 DOWNTO 0);
	sub_wire58    <= data6x(31 DOWNTO 0);
	sub_wire57    <= data7x(31 DOWNTO 0);
	sub_wire56    <= data8x(31 DOWNTO 0);
	sub_wire55    <= data9x(31 DOWNTO 0);
	sub_wire54    <= data10x(31 DOWNTO 0);
	sub_wire53    <= data11x(31 DOWNTO 0);
	sub_wire52    <= data12x(31 DOWNTO 0);
	sub_wire51    <= data13x(31 DOWNTO 0);
	sub_wire50    <= data14x(31 DOWNTO 0);
	sub_wire49    <= data15x(31 DOWNTO 0);
	sub_wire48    <= data16x(31 DOWNTO 0);
	sub_wire47    <= data17x(31 DOWNTO 0);
	sub_wire46    <= data18x(31 DOWNTO 0);
	sub_wire45    <= data19x(31 DOWNTO 0);
	sub_wire44    <= data20x(31 DOWNTO 0);
	sub_wire43    <= data21x(31 DOWNTO 0);
	sub_wire42    <= data22x(31 DOWNTO 0);
	sub_wire41    <= data23x(31 DOWNTO 0);
	sub_wire40    <= data24x(31 DOWNTO 0);
	sub_wire39    <= data25x(31 DOWNTO 0);
	sub_wire38    <= data26x(31 DOWNTO 0);
	sub_wire37    <= data27x(31 DOWNTO 0);
	sub_wire36    <= data28x(31 DOWNTO 0);
	sub_wire35    <= data29x(31 DOWNTO 0);
	sub_wire34    <= data30x(31 DOWNTO 0);
	sub_wire33    <= data31x(31 DOWNTO 0);
	sub_wire32    <= data32x(31 DOWNTO 0);
	sub_wire31    <= data33x(31 DOWNTO 0);
	sub_wire30    <= data34x(31 DOWNTO 0);
	sub_wire29    <= data35x(31 DOWNTO 0);
	sub_wire28    <= data36x(31 DOWNTO 0);
	sub_wire27    <= data37x(31 DOWNTO 0);
	sub_wire26    <= data38x(31 DOWNTO 0);
	sub_wire25    <= data39x(31 DOWNTO 0);
	sub_wire24    <= data40x(31 DOWNTO 0);
	sub_wire23    <= data41x(31 DOWNTO 0);
	sub_wire22    <= data42x(31 DOWNTO 0);
	sub_wire21    <= data43x(31 DOWNTO 0);
	sub_wire20    <= data44x(31 DOWNTO 0);
	sub_wire19    <= data45x(31 DOWNTO 0);
	sub_wire18    <= data46x(31 DOWNTO 0);
	sub_wire17    <= data47x(31 DOWNTO 0);
	sub_wire16    <= data48x(31 DOWNTO 0);
	sub_wire15    <= data49x(31 DOWNTO 0);
	sub_wire14    <= data50x(31 DOWNTO 0);
	sub_wire13    <= data51x(31 DOWNTO 0);
	sub_wire12    <= data52x(31 DOWNTO 0);
	sub_wire11    <= data53x(31 DOWNTO 0);
	sub_wire10    <= data54x(31 DOWNTO 0);
	sub_wire9    <= data55x(31 DOWNTO 0);
	sub_wire8    <= data56x(31 DOWNTO 0);
	sub_wire7    <= data57x(31 DOWNTO 0);
	sub_wire6    <= data58x(31 DOWNTO 0);
	sub_wire5    <= data59x(31 DOWNTO 0);
	sub_wire4    <= data60x(31 DOWNTO 0);
	sub_wire3    <= data61x(31 DOWNTO 0);
	sub_wire2    <= data62x(31 DOWNTO 0);
	sub_wire0    <= data63x(31 DOWNTO 0);
	sub_wire1(63, 0)    <= sub_wire0(0);
	sub_wire1(63, 1)    <= sub_wire0(1);
	sub_wire1(63, 2)    <= sub_wire0(2);
	sub_wire1(63, 3)    <= sub_wire0(3);
	sub_wire1(63, 4)    <= sub_wire0(4);
	sub_wire1(63, 5)    <= sub_wire0(5);
	sub_wire1(63, 6)    <= sub_wire0(6);
	sub_wire1(63, 7)    <= sub_wire0(7);
	sub_wire1(63, 8)    <= sub_wire0(8);
	sub_wire1(63, 9)    <= sub_wire0(9);
	sub_wire1(63, 10)    <= sub_wire0(10);
	sub_wire1(63, 11)    <= sub_wire0(11);
	sub_wire1(63, 12)    <= sub_wire0(12);
	sub_wire1(63, 13)    <= sub_wire0(13);
	sub_wire1(63, 14)    <= sub_wire0(14);
	sub_wire1(63, 15)    <= sub_wire0(15);
	sub_wire1(63, 16)    <= sub_wire0(16);
	sub_wire1(63, 17)    <= sub_wire0(17);
	sub_wire1(63, 18)    <= sub_wire0(18);
	sub_wire1(63, 19)    <= sub_wire0(19);
	sub_wire1(63, 20)    <= sub_wire0(20);
	sub_wire1(63, 21)    <= sub_wire0(21);
	sub_wire1(63, 22)    <= sub_wire0(22);
	sub_wire1(63, 23)    <= sub_wire0(23);
	sub_wire1(63, 24)    <= sub_wire0(24);
	sub_wire1(63, 25)    <= sub_wire0(25);
	sub_wire1(63, 26)    <= sub_wire0(26);
	sub_wire1(63, 27)    <= sub_wire0(27);
	sub_wire1(63, 28)    <= sub_wire0(28);
	sub_wire1(63, 29)    <= sub_wire0(29);
	sub_wire1(63, 30)    <= sub_wire0(30);
	sub_wire1(63, 31)    <= sub_wire0(31);
	sub_wire1(62, 0)    <= sub_wire2(0);
	sub_wire1(62, 1)    <= sub_wire2(1);
	sub_wire1(62, 2)    <= sub_wire2(2);
	sub_wire1(62, 3)    <= sub_wire2(3);
	sub_wire1(62, 4)    <= sub_wire2(4);
	sub_wire1(62, 5)    <= sub_wire2(5);
	sub_wire1(62, 6)    <= sub_wire2(6);
	sub_wire1(62, 7)    <= sub_wire2(7);
	sub_wire1(62, 8)    <= sub_wire2(8);
	sub_wire1(62, 9)    <= sub_wire2(9);
	sub_wire1(62, 10)    <= sub_wire2(10);
	sub_wire1(62, 11)    <= sub_wire2(11);
	sub_wire1(62, 12)    <= sub_wire2(12);
	sub_wire1(62, 13)    <= sub_wire2(13);
	sub_wire1(62, 14)    <= sub_wire2(14);
	sub_wire1(62, 15)    <= sub_wire2(15);
	sub_wire1(62, 16)    <= sub_wire2(16);
	sub_wire1(62, 17)    <= sub_wire2(17);
	sub_wire1(62, 18)    <= sub_wire2(18);
	sub_wire1(62, 19)    <= sub_wire2(19);
	sub_wire1(62, 20)    <= sub_wire2(20);
	sub_wire1(62, 21)    <= sub_wire2(21);
	sub_wire1(62, 22)    <= sub_wire2(22);
	sub_wire1(62, 23)    <= sub_wire2(23);
	sub_wire1(62, 24)    <= sub_wire2(24);
	sub_wire1(62, 25)    <= sub_wire2(25);
	sub_wire1(62, 26)    <= sub_wire2(26);
	sub_wire1(62, 27)    <= sub_wire2(27);
	sub_wire1(62, 28)    <= sub_wire2(28);
	sub_wire1(62, 29)    <= sub_wire2(29);
	sub_wire1(62, 30)    <= sub_wire2(30);
	sub_wire1(62, 31)    <= sub_wire2(31);
	sub_wire1(61, 0)    <= sub_wire3(0);
	sub_wire1(61, 1)    <= sub_wire3(1);
	sub_wire1(61, 2)    <= sub_wire3(2);
	sub_wire1(61, 3)    <= sub_wire3(3);
	sub_wire1(61, 4)    <= sub_wire3(4);
	sub_wire1(61, 5)    <= sub_wire3(5);
	sub_wire1(61, 6)    <= sub_wire3(6);
	sub_wire1(61, 7)    <= sub_wire3(7);
	sub_wire1(61, 8)    <= sub_wire3(8);
	sub_wire1(61, 9)    <= sub_wire3(9);
	sub_wire1(61, 10)    <= sub_wire3(10);
	sub_wire1(61, 11)    <= sub_wire3(11);
	sub_wire1(61, 12)    <= sub_wire3(12);
	sub_wire1(61, 13)    <= sub_wire3(13);
	sub_wire1(61, 14)    <= sub_wire3(14);
	sub_wire1(61, 15)    <= sub_wire3(15);
	sub_wire1(61, 16)    <= sub_wire3(16);
	sub_wire1(61, 17)    <= sub_wire3(17);
	sub_wire1(61, 18)    <= sub_wire3(18);
	sub_wire1(61, 19)    <= sub_wire3(19);
	sub_wire1(61, 20)    <= sub_wire3(20);
	sub_wire1(61, 21)    <= sub_wire3(21);
	sub_wire1(61, 22)    <= sub_wire3(22);
	sub_wire1(61, 23)    <= sub_wire3(23);
	sub_wire1(61, 24)    <= sub_wire3(24);
	sub_wire1(61, 25)    <= sub_wire3(25);
	sub_wire1(61, 26)    <= sub_wire3(26);
	sub_wire1(61, 27)    <= sub_wire3(27);
	sub_wire1(61, 28)    <= sub_wire3(28);
	sub_wire1(61, 29)    <= sub_wire3(29);
	sub_wire1(61, 30)    <= sub_wire3(30);
	sub_wire1(61, 31)    <= sub_wire3(31);
	sub_wire1(60, 0)    <= sub_wire4(0);
	sub_wire1(60, 1)    <= sub_wire4(1);
	sub_wire1(60, 2)    <= sub_wire4(2);
	sub_wire1(60, 3)    <= sub_wire4(3);
	sub_wire1(60, 4)    <= sub_wire4(4);
	sub_wire1(60, 5)    <= sub_wire4(5);
	sub_wire1(60, 6)    <= sub_wire4(6);
	sub_wire1(60, 7)    <= sub_wire4(7);
	sub_wire1(60, 8)    <= sub_wire4(8);
	sub_wire1(60, 9)    <= sub_wire4(9);
	sub_wire1(60, 10)    <= sub_wire4(10);
	sub_wire1(60, 11)    <= sub_wire4(11);
	sub_wire1(60, 12)    <= sub_wire4(12);
	sub_wire1(60, 13)    <= sub_wire4(13);
	sub_wire1(60, 14)    <= sub_wire4(14);
	sub_wire1(60, 15)    <= sub_wire4(15);
	sub_wire1(60, 16)    <= sub_wire4(16);
	sub_wire1(60, 17)    <= sub_wire4(17);
	sub_wire1(60, 18)    <= sub_wire4(18);
	sub_wire1(60, 19)    <= sub_wire4(19);
	sub_wire1(60, 20)    <= sub_wire4(20);
	sub_wire1(60, 21)    <= sub_wire4(21);
	sub_wire1(60, 22)    <= sub_wire4(22);
	sub_wire1(60, 23)    <= sub_wire4(23);
	sub_wire1(60, 24)    <= sub_wire4(24);
	sub_wire1(60, 25)    <= sub_wire4(25);
	sub_wire1(60, 26)    <= sub_wire4(26);
	sub_wire1(60, 27)    <= sub_wire4(27);
	sub_wire1(60, 28)    <= sub_wire4(28);
	sub_wire1(60, 29)    <= sub_wire4(29);
	sub_wire1(60, 30)    <= sub_wire4(30);
	sub_wire1(60, 31)    <= sub_wire4(31);
	sub_wire1(59, 0)    <= sub_wire5(0);
	sub_wire1(59, 1)    <= sub_wire5(1);
	sub_wire1(59, 2)    <= sub_wire5(2);
	sub_wire1(59, 3)    <= sub_wire5(3);
	sub_wire1(59, 4)    <= sub_wire5(4);
	sub_wire1(59, 5)    <= sub_wire5(5);
	sub_wire1(59, 6)    <= sub_wire5(6);
	sub_wire1(59, 7)    <= sub_wire5(7);
	sub_wire1(59, 8)    <= sub_wire5(8);
	sub_wire1(59, 9)    <= sub_wire5(9);
	sub_wire1(59, 10)    <= sub_wire5(10);
	sub_wire1(59, 11)    <= sub_wire5(11);
	sub_wire1(59, 12)    <= sub_wire5(12);
	sub_wire1(59, 13)    <= sub_wire5(13);
	sub_wire1(59, 14)    <= sub_wire5(14);
	sub_wire1(59, 15)    <= sub_wire5(15);
	sub_wire1(59, 16)    <= sub_wire5(16);
	sub_wire1(59, 17)    <= sub_wire5(17);
	sub_wire1(59, 18)    <= sub_wire5(18);
	sub_wire1(59, 19)    <= sub_wire5(19);
	sub_wire1(59, 20)    <= sub_wire5(20);
	sub_wire1(59, 21)    <= sub_wire5(21);
	sub_wire1(59, 22)    <= sub_wire5(22);
	sub_wire1(59, 23)    <= sub_wire5(23);
	sub_wire1(59, 24)    <= sub_wire5(24);
	sub_wire1(59, 25)    <= sub_wire5(25);
	sub_wire1(59, 26)    <= sub_wire5(26);
	sub_wire1(59, 27)    <= sub_wire5(27);
	sub_wire1(59, 28)    <= sub_wire5(28);
	sub_wire1(59, 29)    <= sub_wire5(29);
	sub_wire1(59, 30)    <= sub_wire5(30);
	sub_wire1(59, 31)    <= sub_wire5(31);
	sub_wire1(58, 0)    <= sub_wire6(0);
	sub_wire1(58, 1)    <= sub_wire6(1);
	sub_wire1(58, 2)    <= sub_wire6(2);
	sub_wire1(58, 3)    <= sub_wire6(3);
	sub_wire1(58, 4)    <= sub_wire6(4);
	sub_wire1(58, 5)    <= sub_wire6(5);
	sub_wire1(58, 6)    <= sub_wire6(6);
	sub_wire1(58, 7)    <= sub_wire6(7);
	sub_wire1(58, 8)    <= sub_wire6(8);
	sub_wire1(58, 9)    <= sub_wire6(9);
	sub_wire1(58, 10)    <= sub_wire6(10);
	sub_wire1(58, 11)    <= sub_wire6(11);
	sub_wire1(58, 12)    <= sub_wire6(12);
	sub_wire1(58, 13)    <= sub_wire6(13);
	sub_wire1(58, 14)    <= sub_wire6(14);
	sub_wire1(58, 15)    <= sub_wire6(15);
	sub_wire1(58, 16)    <= sub_wire6(16);
	sub_wire1(58, 17)    <= sub_wire6(17);
	sub_wire1(58, 18)    <= sub_wire6(18);
	sub_wire1(58, 19)    <= sub_wire6(19);
	sub_wire1(58, 20)    <= sub_wire6(20);
	sub_wire1(58, 21)    <= sub_wire6(21);
	sub_wire1(58, 22)    <= sub_wire6(22);
	sub_wire1(58, 23)    <= sub_wire6(23);
	sub_wire1(58, 24)    <= sub_wire6(24);
	sub_wire1(58, 25)    <= sub_wire6(25);
	sub_wire1(58, 26)    <= sub_wire6(26);
	sub_wire1(58, 27)    <= sub_wire6(27);
	sub_wire1(58, 28)    <= sub_wire6(28);
	sub_wire1(58, 29)    <= sub_wire6(29);
	sub_wire1(58, 30)    <= sub_wire6(30);
	sub_wire1(58, 31)    <= sub_wire6(31);
	sub_wire1(57, 0)    <= sub_wire7(0);
	sub_wire1(57, 1)    <= sub_wire7(1);
	sub_wire1(57, 2)    <= sub_wire7(2);
	sub_wire1(57, 3)    <= sub_wire7(3);
	sub_wire1(57, 4)    <= sub_wire7(4);
	sub_wire1(57, 5)    <= sub_wire7(5);
	sub_wire1(57, 6)    <= sub_wire7(6);
	sub_wire1(57, 7)    <= sub_wire7(7);
	sub_wire1(57, 8)    <= sub_wire7(8);
	sub_wire1(57, 9)    <= sub_wire7(9);
	sub_wire1(57, 10)    <= sub_wire7(10);
	sub_wire1(57, 11)    <= sub_wire7(11);
	sub_wire1(57, 12)    <= sub_wire7(12);
	sub_wire1(57, 13)    <= sub_wire7(13);
	sub_wire1(57, 14)    <= sub_wire7(14);
	sub_wire1(57, 15)    <= sub_wire7(15);
	sub_wire1(57, 16)    <= sub_wire7(16);
	sub_wire1(57, 17)    <= sub_wire7(17);
	sub_wire1(57, 18)    <= sub_wire7(18);
	sub_wire1(57, 19)    <= sub_wire7(19);
	sub_wire1(57, 20)    <= sub_wire7(20);
	sub_wire1(57, 21)    <= sub_wire7(21);
	sub_wire1(57, 22)    <= sub_wire7(22);
	sub_wire1(57, 23)    <= sub_wire7(23);
	sub_wire1(57, 24)    <= sub_wire7(24);
	sub_wire1(57, 25)    <= sub_wire7(25);
	sub_wire1(57, 26)    <= sub_wire7(26);
	sub_wire1(57, 27)    <= sub_wire7(27);
	sub_wire1(57, 28)    <= sub_wire7(28);
	sub_wire1(57, 29)    <= sub_wire7(29);
	sub_wire1(57, 30)    <= sub_wire7(30);
	sub_wire1(57, 31)    <= sub_wire7(31);
	sub_wire1(56, 0)    <= sub_wire8(0);
	sub_wire1(56, 1)    <= sub_wire8(1);
	sub_wire1(56, 2)    <= sub_wire8(2);
	sub_wire1(56, 3)    <= sub_wire8(3);
	sub_wire1(56, 4)    <= sub_wire8(4);
	sub_wire1(56, 5)    <= sub_wire8(5);
	sub_wire1(56, 6)    <= sub_wire8(6);
	sub_wire1(56, 7)    <= sub_wire8(7);
	sub_wire1(56, 8)    <= sub_wire8(8);
	sub_wire1(56, 9)    <= sub_wire8(9);
	sub_wire1(56, 10)    <= sub_wire8(10);
	sub_wire1(56, 11)    <= sub_wire8(11);
	sub_wire1(56, 12)    <= sub_wire8(12);
	sub_wire1(56, 13)    <= sub_wire8(13);
	sub_wire1(56, 14)    <= sub_wire8(14);
	sub_wire1(56, 15)    <= sub_wire8(15);
	sub_wire1(56, 16)    <= sub_wire8(16);
	sub_wire1(56, 17)    <= sub_wire8(17);
	sub_wire1(56, 18)    <= sub_wire8(18);
	sub_wire1(56, 19)    <= sub_wire8(19);
	sub_wire1(56, 20)    <= sub_wire8(20);
	sub_wire1(56, 21)    <= sub_wire8(21);
	sub_wire1(56, 22)    <= sub_wire8(22);
	sub_wire1(56, 23)    <= sub_wire8(23);
	sub_wire1(56, 24)    <= sub_wire8(24);
	sub_wire1(56, 25)    <= sub_wire8(25);
	sub_wire1(56, 26)    <= sub_wire8(26);
	sub_wire1(56, 27)    <= sub_wire8(27);
	sub_wire1(56, 28)    <= sub_wire8(28);
	sub_wire1(56, 29)    <= sub_wire8(29);
	sub_wire1(56, 30)    <= sub_wire8(30);
	sub_wire1(56, 31)    <= sub_wire8(31);
	sub_wire1(55, 0)    <= sub_wire9(0);
	sub_wire1(55, 1)    <= sub_wire9(1);
	sub_wire1(55, 2)    <= sub_wire9(2);
	sub_wire1(55, 3)    <= sub_wire9(3);
	sub_wire1(55, 4)    <= sub_wire9(4);
	sub_wire1(55, 5)    <= sub_wire9(5);
	sub_wire1(55, 6)    <= sub_wire9(6);
	sub_wire1(55, 7)    <= sub_wire9(7);
	sub_wire1(55, 8)    <= sub_wire9(8);
	sub_wire1(55, 9)    <= sub_wire9(9);
	sub_wire1(55, 10)    <= sub_wire9(10);
	sub_wire1(55, 11)    <= sub_wire9(11);
	sub_wire1(55, 12)    <= sub_wire9(12);
	sub_wire1(55, 13)    <= sub_wire9(13);
	sub_wire1(55, 14)    <= sub_wire9(14);
	sub_wire1(55, 15)    <= sub_wire9(15);
	sub_wire1(55, 16)    <= sub_wire9(16);
	sub_wire1(55, 17)    <= sub_wire9(17);
	sub_wire1(55, 18)    <= sub_wire9(18);
	sub_wire1(55, 19)    <= sub_wire9(19);
	sub_wire1(55, 20)    <= sub_wire9(20);
	sub_wire1(55, 21)    <= sub_wire9(21);
	sub_wire1(55, 22)    <= sub_wire9(22);
	sub_wire1(55, 23)    <= sub_wire9(23);
	sub_wire1(55, 24)    <= sub_wire9(24);
	sub_wire1(55, 25)    <= sub_wire9(25);
	sub_wire1(55, 26)    <= sub_wire9(26);
	sub_wire1(55, 27)    <= sub_wire9(27);
	sub_wire1(55, 28)    <= sub_wire9(28);
	sub_wire1(55, 29)    <= sub_wire9(29);
	sub_wire1(55, 30)    <= sub_wire9(30);
	sub_wire1(55, 31)    <= sub_wire9(31);
	sub_wire1(54, 0)    <= sub_wire10(0);
	sub_wire1(54, 1)    <= sub_wire10(1);
	sub_wire1(54, 2)    <= sub_wire10(2);
	sub_wire1(54, 3)    <= sub_wire10(3);
	sub_wire1(54, 4)    <= sub_wire10(4);
	sub_wire1(54, 5)    <= sub_wire10(5);
	sub_wire1(54, 6)    <= sub_wire10(6);
	sub_wire1(54, 7)    <= sub_wire10(7);
	sub_wire1(54, 8)    <= sub_wire10(8);
	sub_wire1(54, 9)    <= sub_wire10(9);
	sub_wire1(54, 10)    <= sub_wire10(10);
	sub_wire1(54, 11)    <= sub_wire10(11);
	sub_wire1(54, 12)    <= sub_wire10(12);
	sub_wire1(54, 13)    <= sub_wire10(13);
	sub_wire1(54, 14)    <= sub_wire10(14);
	sub_wire1(54, 15)    <= sub_wire10(15);
	sub_wire1(54, 16)    <= sub_wire10(16);
	sub_wire1(54, 17)    <= sub_wire10(17);
	sub_wire1(54, 18)    <= sub_wire10(18);
	sub_wire1(54, 19)    <= sub_wire10(19);
	sub_wire1(54, 20)    <= sub_wire10(20);
	sub_wire1(54, 21)    <= sub_wire10(21);
	sub_wire1(54, 22)    <= sub_wire10(22);
	sub_wire1(54, 23)    <= sub_wire10(23);
	sub_wire1(54, 24)    <= sub_wire10(24);
	sub_wire1(54, 25)    <= sub_wire10(25);
	sub_wire1(54, 26)    <= sub_wire10(26);
	sub_wire1(54, 27)    <= sub_wire10(27);
	sub_wire1(54, 28)    <= sub_wire10(28);
	sub_wire1(54, 29)    <= sub_wire10(29);
	sub_wire1(54, 30)    <= sub_wire10(30);
	sub_wire1(54, 31)    <= sub_wire10(31);
	sub_wire1(53, 0)    <= sub_wire11(0);
	sub_wire1(53, 1)    <= sub_wire11(1);
	sub_wire1(53, 2)    <= sub_wire11(2);
	sub_wire1(53, 3)    <= sub_wire11(3);
	sub_wire1(53, 4)    <= sub_wire11(4);
	sub_wire1(53, 5)    <= sub_wire11(5);
	sub_wire1(53, 6)    <= sub_wire11(6);
	sub_wire1(53, 7)    <= sub_wire11(7);
	sub_wire1(53, 8)    <= sub_wire11(8);
	sub_wire1(53, 9)    <= sub_wire11(9);
	sub_wire1(53, 10)    <= sub_wire11(10);
	sub_wire1(53, 11)    <= sub_wire11(11);
	sub_wire1(53, 12)    <= sub_wire11(12);
	sub_wire1(53, 13)    <= sub_wire11(13);
	sub_wire1(53, 14)    <= sub_wire11(14);
	sub_wire1(53, 15)    <= sub_wire11(15);
	sub_wire1(53, 16)    <= sub_wire11(16);
	sub_wire1(53, 17)    <= sub_wire11(17);
	sub_wire1(53, 18)    <= sub_wire11(18);
	sub_wire1(53, 19)    <= sub_wire11(19);
	sub_wire1(53, 20)    <= sub_wire11(20);
	sub_wire1(53, 21)    <= sub_wire11(21);
	sub_wire1(53, 22)    <= sub_wire11(22);
	sub_wire1(53, 23)    <= sub_wire11(23);
	sub_wire1(53, 24)    <= sub_wire11(24);
	sub_wire1(53, 25)    <= sub_wire11(25);
	sub_wire1(53, 26)    <= sub_wire11(26);
	sub_wire1(53, 27)    <= sub_wire11(27);
	sub_wire1(53, 28)    <= sub_wire11(28);
	sub_wire1(53, 29)    <= sub_wire11(29);
	sub_wire1(53, 30)    <= sub_wire11(30);
	sub_wire1(53, 31)    <= sub_wire11(31);
	sub_wire1(52, 0)    <= sub_wire12(0);
	sub_wire1(52, 1)    <= sub_wire12(1);
	sub_wire1(52, 2)    <= sub_wire12(2);
	sub_wire1(52, 3)    <= sub_wire12(3);
	sub_wire1(52, 4)    <= sub_wire12(4);
	sub_wire1(52, 5)    <= sub_wire12(5);
	sub_wire1(52, 6)    <= sub_wire12(6);
	sub_wire1(52, 7)    <= sub_wire12(7);
	sub_wire1(52, 8)    <= sub_wire12(8);
	sub_wire1(52, 9)    <= sub_wire12(9);
	sub_wire1(52, 10)    <= sub_wire12(10);
	sub_wire1(52, 11)    <= sub_wire12(11);
	sub_wire1(52, 12)    <= sub_wire12(12);
	sub_wire1(52, 13)    <= sub_wire12(13);
	sub_wire1(52, 14)    <= sub_wire12(14);
	sub_wire1(52, 15)    <= sub_wire12(15);
	sub_wire1(52, 16)    <= sub_wire12(16);
	sub_wire1(52, 17)    <= sub_wire12(17);
	sub_wire1(52, 18)    <= sub_wire12(18);
	sub_wire1(52, 19)    <= sub_wire12(19);
	sub_wire1(52, 20)    <= sub_wire12(20);
	sub_wire1(52, 21)    <= sub_wire12(21);
	sub_wire1(52, 22)    <= sub_wire12(22);
	sub_wire1(52, 23)    <= sub_wire12(23);
	sub_wire1(52, 24)    <= sub_wire12(24);
	sub_wire1(52, 25)    <= sub_wire12(25);
	sub_wire1(52, 26)    <= sub_wire12(26);
	sub_wire1(52, 27)    <= sub_wire12(27);
	sub_wire1(52, 28)    <= sub_wire12(28);
	sub_wire1(52, 29)    <= sub_wire12(29);
	sub_wire1(52, 30)    <= sub_wire12(30);
	sub_wire1(52, 31)    <= sub_wire12(31);
	sub_wire1(51, 0)    <= sub_wire13(0);
	sub_wire1(51, 1)    <= sub_wire13(1);
	sub_wire1(51, 2)    <= sub_wire13(2);
	sub_wire1(51, 3)    <= sub_wire13(3);
	sub_wire1(51, 4)    <= sub_wire13(4);
	sub_wire1(51, 5)    <= sub_wire13(5);
	sub_wire1(51, 6)    <= sub_wire13(6);
	sub_wire1(51, 7)    <= sub_wire13(7);
	sub_wire1(51, 8)    <= sub_wire13(8);
	sub_wire1(51, 9)    <= sub_wire13(9);
	sub_wire1(51, 10)    <= sub_wire13(10);
	sub_wire1(51, 11)    <= sub_wire13(11);
	sub_wire1(51, 12)    <= sub_wire13(12);
	sub_wire1(51, 13)    <= sub_wire13(13);
	sub_wire1(51, 14)    <= sub_wire13(14);
	sub_wire1(51, 15)    <= sub_wire13(15);
	sub_wire1(51, 16)    <= sub_wire13(16);
	sub_wire1(51, 17)    <= sub_wire13(17);
	sub_wire1(51, 18)    <= sub_wire13(18);
	sub_wire1(51, 19)    <= sub_wire13(19);
	sub_wire1(51, 20)    <= sub_wire13(20);
	sub_wire1(51, 21)    <= sub_wire13(21);
	sub_wire1(51, 22)    <= sub_wire13(22);
	sub_wire1(51, 23)    <= sub_wire13(23);
	sub_wire1(51, 24)    <= sub_wire13(24);
	sub_wire1(51, 25)    <= sub_wire13(25);
	sub_wire1(51, 26)    <= sub_wire13(26);
	sub_wire1(51, 27)    <= sub_wire13(27);
	sub_wire1(51, 28)    <= sub_wire13(28);
	sub_wire1(51, 29)    <= sub_wire13(29);
	sub_wire1(51, 30)    <= sub_wire13(30);
	sub_wire1(51, 31)    <= sub_wire13(31);
	sub_wire1(50, 0)    <= sub_wire14(0);
	sub_wire1(50, 1)    <= sub_wire14(1);
	sub_wire1(50, 2)    <= sub_wire14(2);
	sub_wire1(50, 3)    <= sub_wire14(3);
	sub_wire1(50, 4)    <= sub_wire14(4);
	sub_wire1(50, 5)    <= sub_wire14(5);
	sub_wire1(50, 6)    <= sub_wire14(6);
	sub_wire1(50, 7)    <= sub_wire14(7);
	sub_wire1(50, 8)    <= sub_wire14(8);
	sub_wire1(50, 9)    <= sub_wire14(9);
	sub_wire1(50, 10)    <= sub_wire14(10);
	sub_wire1(50, 11)    <= sub_wire14(11);
	sub_wire1(50, 12)    <= sub_wire14(12);
	sub_wire1(50, 13)    <= sub_wire14(13);
	sub_wire1(50, 14)    <= sub_wire14(14);
	sub_wire1(50, 15)    <= sub_wire14(15);
	sub_wire1(50, 16)    <= sub_wire14(16);
	sub_wire1(50, 17)    <= sub_wire14(17);
	sub_wire1(50, 18)    <= sub_wire14(18);
	sub_wire1(50, 19)    <= sub_wire14(19);
	sub_wire1(50, 20)    <= sub_wire14(20);
	sub_wire1(50, 21)    <= sub_wire14(21);
	sub_wire1(50, 22)    <= sub_wire14(22);
	sub_wire1(50, 23)    <= sub_wire14(23);
	sub_wire1(50, 24)    <= sub_wire14(24);
	sub_wire1(50, 25)    <= sub_wire14(25);
	sub_wire1(50, 26)    <= sub_wire14(26);
	sub_wire1(50, 27)    <= sub_wire14(27);
	sub_wire1(50, 28)    <= sub_wire14(28);
	sub_wire1(50, 29)    <= sub_wire14(29);
	sub_wire1(50, 30)    <= sub_wire14(30);
	sub_wire1(50, 31)    <= sub_wire14(31);
	sub_wire1(49, 0)    <= sub_wire15(0);
	sub_wire1(49, 1)    <= sub_wire15(1);
	sub_wire1(49, 2)    <= sub_wire15(2);
	sub_wire1(49, 3)    <= sub_wire15(3);
	sub_wire1(49, 4)    <= sub_wire15(4);
	sub_wire1(49, 5)    <= sub_wire15(5);
	sub_wire1(49, 6)    <= sub_wire15(6);
	sub_wire1(49, 7)    <= sub_wire15(7);
	sub_wire1(49, 8)    <= sub_wire15(8);
	sub_wire1(49, 9)    <= sub_wire15(9);
	sub_wire1(49, 10)    <= sub_wire15(10);
	sub_wire1(49, 11)    <= sub_wire15(11);
	sub_wire1(49, 12)    <= sub_wire15(12);
	sub_wire1(49, 13)    <= sub_wire15(13);
	sub_wire1(49, 14)    <= sub_wire15(14);
	sub_wire1(49, 15)    <= sub_wire15(15);
	sub_wire1(49, 16)    <= sub_wire15(16);
	sub_wire1(49, 17)    <= sub_wire15(17);
	sub_wire1(49, 18)    <= sub_wire15(18);
	sub_wire1(49, 19)    <= sub_wire15(19);
	sub_wire1(49, 20)    <= sub_wire15(20);
	sub_wire1(49, 21)    <= sub_wire15(21);
	sub_wire1(49, 22)    <= sub_wire15(22);
	sub_wire1(49, 23)    <= sub_wire15(23);
	sub_wire1(49, 24)    <= sub_wire15(24);
	sub_wire1(49, 25)    <= sub_wire15(25);
	sub_wire1(49, 26)    <= sub_wire15(26);
	sub_wire1(49, 27)    <= sub_wire15(27);
	sub_wire1(49, 28)    <= sub_wire15(28);
	sub_wire1(49, 29)    <= sub_wire15(29);
	sub_wire1(49, 30)    <= sub_wire15(30);
	sub_wire1(49, 31)    <= sub_wire15(31);
	sub_wire1(48, 0)    <= sub_wire16(0);
	sub_wire1(48, 1)    <= sub_wire16(1);
	sub_wire1(48, 2)    <= sub_wire16(2);
	sub_wire1(48, 3)    <= sub_wire16(3);
	sub_wire1(48, 4)    <= sub_wire16(4);
	sub_wire1(48, 5)    <= sub_wire16(5);
	sub_wire1(48, 6)    <= sub_wire16(6);
	sub_wire1(48, 7)    <= sub_wire16(7);
	sub_wire1(48, 8)    <= sub_wire16(8);
	sub_wire1(48, 9)    <= sub_wire16(9);
	sub_wire1(48, 10)    <= sub_wire16(10);
	sub_wire1(48, 11)    <= sub_wire16(11);
	sub_wire1(48, 12)    <= sub_wire16(12);
	sub_wire1(48, 13)    <= sub_wire16(13);
	sub_wire1(48, 14)    <= sub_wire16(14);
	sub_wire1(48, 15)    <= sub_wire16(15);
	sub_wire1(48, 16)    <= sub_wire16(16);
	sub_wire1(48, 17)    <= sub_wire16(17);
	sub_wire1(48, 18)    <= sub_wire16(18);
	sub_wire1(48, 19)    <= sub_wire16(19);
	sub_wire1(48, 20)    <= sub_wire16(20);
	sub_wire1(48, 21)    <= sub_wire16(21);
	sub_wire1(48, 22)    <= sub_wire16(22);
	sub_wire1(48, 23)    <= sub_wire16(23);
	sub_wire1(48, 24)    <= sub_wire16(24);
	sub_wire1(48, 25)    <= sub_wire16(25);
	sub_wire1(48, 26)    <= sub_wire16(26);
	sub_wire1(48, 27)    <= sub_wire16(27);
	sub_wire1(48, 28)    <= sub_wire16(28);
	sub_wire1(48, 29)    <= sub_wire16(29);
	sub_wire1(48, 30)    <= sub_wire16(30);
	sub_wire1(48, 31)    <= sub_wire16(31);
	sub_wire1(47, 0)    <= sub_wire17(0);
	sub_wire1(47, 1)    <= sub_wire17(1);
	sub_wire1(47, 2)    <= sub_wire17(2);
	sub_wire1(47, 3)    <= sub_wire17(3);
	sub_wire1(47, 4)    <= sub_wire17(4);
	sub_wire1(47, 5)    <= sub_wire17(5);
	sub_wire1(47, 6)    <= sub_wire17(6);
	sub_wire1(47, 7)    <= sub_wire17(7);
	sub_wire1(47, 8)    <= sub_wire17(8);
	sub_wire1(47, 9)    <= sub_wire17(9);
	sub_wire1(47, 10)    <= sub_wire17(10);
	sub_wire1(47, 11)    <= sub_wire17(11);
	sub_wire1(47, 12)    <= sub_wire17(12);
	sub_wire1(47, 13)    <= sub_wire17(13);
	sub_wire1(47, 14)    <= sub_wire17(14);
	sub_wire1(47, 15)    <= sub_wire17(15);
	sub_wire1(47, 16)    <= sub_wire17(16);
	sub_wire1(47, 17)    <= sub_wire17(17);
	sub_wire1(47, 18)    <= sub_wire17(18);
	sub_wire1(47, 19)    <= sub_wire17(19);
	sub_wire1(47, 20)    <= sub_wire17(20);
	sub_wire1(47, 21)    <= sub_wire17(21);
	sub_wire1(47, 22)    <= sub_wire17(22);
	sub_wire1(47, 23)    <= sub_wire17(23);
	sub_wire1(47, 24)    <= sub_wire17(24);
	sub_wire1(47, 25)    <= sub_wire17(25);
	sub_wire1(47, 26)    <= sub_wire17(26);
	sub_wire1(47, 27)    <= sub_wire17(27);
	sub_wire1(47, 28)    <= sub_wire17(28);
	sub_wire1(47, 29)    <= sub_wire17(29);
	sub_wire1(47, 30)    <= sub_wire17(30);
	sub_wire1(47, 31)    <= sub_wire17(31);
	sub_wire1(46, 0)    <= sub_wire18(0);
	sub_wire1(46, 1)    <= sub_wire18(1);
	sub_wire1(46, 2)    <= sub_wire18(2);
	sub_wire1(46, 3)    <= sub_wire18(3);
	sub_wire1(46, 4)    <= sub_wire18(4);
	sub_wire1(46, 5)    <= sub_wire18(5);
	sub_wire1(46, 6)    <= sub_wire18(6);
	sub_wire1(46, 7)    <= sub_wire18(7);
	sub_wire1(46, 8)    <= sub_wire18(8);
	sub_wire1(46, 9)    <= sub_wire18(9);
	sub_wire1(46, 10)    <= sub_wire18(10);
	sub_wire1(46, 11)    <= sub_wire18(11);
	sub_wire1(46, 12)    <= sub_wire18(12);
	sub_wire1(46, 13)    <= sub_wire18(13);
	sub_wire1(46, 14)    <= sub_wire18(14);
	sub_wire1(46, 15)    <= sub_wire18(15);
	sub_wire1(46, 16)    <= sub_wire18(16);
	sub_wire1(46, 17)    <= sub_wire18(17);
	sub_wire1(46, 18)    <= sub_wire18(18);
	sub_wire1(46, 19)    <= sub_wire18(19);
	sub_wire1(46, 20)    <= sub_wire18(20);
	sub_wire1(46, 21)    <= sub_wire18(21);
	sub_wire1(46, 22)    <= sub_wire18(22);
	sub_wire1(46, 23)    <= sub_wire18(23);
	sub_wire1(46, 24)    <= sub_wire18(24);
	sub_wire1(46, 25)    <= sub_wire18(25);
	sub_wire1(46, 26)    <= sub_wire18(26);
	sub_wire1(46, 27)    <= sub_wire18(27);
	sub_wire1(46, 28)    <= sub_wire18(28);
	sub_wire1(46, 29)    <= sub_wire18(29);
	sub_wire1(46, 30)    <= sub_wire18(30);
	sub_wire1(46, 31)    <= sub_wire18(31);
	sub_wire1(45, 0)    <= sub_wire19(0);
	sub_wire1(45, 1)    <= sub_wire19(1);
	sub_wire1(45, 2)    <= sub_wire19(2);
	sub_wire1(45, 3)    <= sub_wire19(3);
	sub_wire1(45, 4)    <= sub_wire19(4);
	sub_wire1(45, 5)    <= sub_wire19(5);
	sub_wire1(45, 6)    <= sub_wire19(6);
	sub_wire1(45, 7)    <= sub_wire19(7);
	sub_wire1(45, 8)    <= sub_wire19(8);
	sub_wire1(45, 9)    <= sub_wire19(9);
	sub_wire1(45, 10)    <= sub_wire19(10);
	sub_wire1(45, 11)    <= sub_wire19(11);
	sub_wire1(45, 12)    <= sub_wire19(12);
	sub_wire1(45, 13)    <= sub_wire19(13);
	sub_wire1(45, 14)    <= sub_wire19(14);
	sub_wire1(45, 15)    <= sub_wire19(15);
	sub_wire1(45, 16)    <= sub_wire19(16);
	sub_wire1(45, 17)    <= sub_wire19(17);
	sub_wire1(45, 18)    <= sub_wire19(18);
	sub_wire1(45, 19)    <= sub_wire19(19);
	sub_wire1(45, 20)    <= sub_wire19(20);
	sub_wire1(45, 21)    <= sub_wire19(21);
	sub_wire1(45, 22)    <= sub_wire19(22);
	sub_wire1(45, 23)    <= sub_wire19(23);
	sub_wire1(45, 24)    <= sub_wire19(24);
	sub_wire1(45, 25)    <= sub_wire19(25);
	sub_wire1(45, 26)    <= sub_wire19(26);
	sub_wire1(45, 27)    <= sub_wire19(27);
	sub_wire1(45, 28)    <= sub_wire19(28);
	sub_wire1(45, 29)    <= sub_wire19(29);
	sub_wire1(45, 30)    <= sub_wire19(30);
	sub_wire1(45, 31)    <= sub_wire19(31);
	sub_wire1(44, 0)    <= sub_wire20(0);
	sub_wire1(44, 1)    <= sub_wire20(1);
	sub_wire1(44, 2)    <= sub_wire20(2);
	sub_wire1(44, 3)    <= sub_wire20(3);
	sub_wire1(44, 4)    <= sub_wire20(4);
	sub_wire1(44, 5)    <= sub_wire20(5);
	sub_wire1(44, 6)    <= sub_wire20(6);
	sub_wire1(44, 7)    <= sub_wire20(7);
	sub_wire1(44, 8)    <= sub_wire20(8);
	sub_wire1(44, 9)    <= sub_wire20(9);
	sub_wire1(44, 10)    <= sub_wire20(10);
	sub_wire1(44, 11)    <= sub_wire20(11);
	sub_wire1(44, 12)    <= sub_wire20(12);
	sub_wire1(44, 13)    <= sub_wire20(13);
	sub_wire1(44, 14)    <= sub_wire20(14);
	sub_wire1(44, 15)    <= sub_wire20(15);
	sub_wire1(44, 16)    <= sub_wire20(16);
	sub_wire1(44, 17)    <= sub_wire20(17);
	sub_wire1(44, 18)    <= sub_wire20(18);
	sub_wire1(44, 19)    <= sub_wire20(19);
	sub_wire1(44, 20)    <= sub_wire20(20);
	sub_wire1(44, 21)    <= sub_wire20(21);
	sub_wire1(44, 22)    <= sub_wire20(22);
	sub_wire1(44, 23)    <= sub_wire20(23);
	sub_wire1(44, 24)    <= sub_wire20(24);
	sub_wire1(44, 25)    <= sub_wire20(25);
	sub_wire1(44, 26)    <= sub_wire20(26);
	sub_wire1(44, 27)    <= sub_wire20(27);
	sub_wire1(44, 28)    <= sub_wire20(28);
	sub_wire1(44, 29)    <= sub_wire20(29);
	sub_wire1(44, 30)    <= sub_wire20(30);
	sub_wire1(44, 31)    <= sub_wire20(31);
	sub_wire1(43, 0)    <= sub_wire21(0);
	sub_wire1(43, 1)    <= sub_wire21(1);
	sub_wire1(43, 2)    <= sub_wire21(2);
	sub_wire1(43, 3)    <= sub_wire21(3);
	sub_wire1(43, 4)    <= sub_wire21(4);
	sub_wire1(43, 5)    <= sub_wire21(5);
	sub_wire1(43, 6)    <= sub_wire21(6);
	sub_wire1(43, 7)    <= sub_wire21(7);
	sub_wire1(43, 8)    <= sub_wire21(8);
	sub_wire1(43, 9)    <= sub_wire21(9);
	sub_wire1(43, 10)    <= sub_wire21(10);
	sub_wire1(43, 11)    <= sub_wire21(11);
	sub_wire1(43, 12)    <= sub_wire21(12);
	sub_wire1(43, 13)    <= sub_wire21(13);
	sub_wire1(43, 14)    <= sub_wire21(14);
	sub_wire1(43, 15)    <= sub_wire21(15);
	sub_wire1(43, 16)    <= sub_wire21(16);
	sub_wire1(43, 17)    <= sub_wire21(17);
	sub_wire1(43, 18)    <= sub_wire21(18);
	sub_wire1(43, 19)    <= sub_wire21(19);
	sub_wire1(43, 20)    <= sub_wire21(20);
	sub_wire1(43, 21)    <= sub_wire21(21);
	sub_wire1(43, 22)    <= sub_wire21(22);
	sub_wire1(43, 23)    <= sub_wire21(23);
	sub_wire1(43, 24)    <= sub_wire21(24);
	sub_wire1(43, 25)    <= sub_wire21(25);
	sub_wire1(43, 26)    <= sub_wire21(26);
	sub_wire1(43, 27)    <= sub_wire21(27);
	sub_wire1(43, 28)    <= sub_wire21(28);
	sub_wire1(43, 29)    <= sub_wire21(29);
	sub_wire1(43, 30)    <= sub_wire21(30);
	sub_wire1(43, 31)    <= sub_wire21(31);
	sub_wire1(42, 0)    <= sub_wire22(0);
	sub_wire1(42, 1)    <= sub_wire22(1);
	sub_wire1(42, 2)    <= sub_wire22(2);
	sub_wire1(42, 3)    <= sub_wire22(3);
	sub_wire1(42, 4)    <= sub_wire22(4);
	sub_wire1(42, 5)    <= sub_wire22(5);
	sub_wire1(42, 6)    <= sub_wire22(6);
	sub_wire1(42, 7)    <= sub_wire22(7);
	sub_wire1(42, 8)    <= sub_wire22(8);
	sub_wire1(42, 9)    <= sub_wire22(9);
	sub_wire1(42, 10)    <= sub_wire22(10);
	sub_wire1(42, 11)    <= sub_wire22(11);
	sub_wire1(42, 12)    <= sub_wire22(12);
	sub_wire1(42, 13)    <= sub_wire22(13);
	sub_wire1(42, 14)    <= sub_wire22(14);
	sub_wire1(42, 15)    <= sub_wire22(15);
	sub_wire1(42, 16)    <= sub_wire22(16);
	sub_wire1(42, 17)    <= sub_wire22(17);
	sub_wire1(42, 18)    <= sub_wire22(18);
	sub_wire1(42, 19)    <= sub_wire22(19);
	sub_wire1(42, 20)    <= sub_wire22(20);
	sub_wire1(42, 21)    <= sub_wire22(21);
	sub_wire1(42, 22)    <= sub_wire22(22);
	sub_wire1(42, 23)    <= sub_wire22(23);
	sub_wire1(42, 24)    <= sub_wire22(24);
	sub_wire1(42, 25)    <= sub_wire22(25);
	sub_wire1(42, 26)    <= sub_wire22(26);
	sub_wire1(42, 27)    <= sub_wire22(27);
	sub_wire1(42, 28)    <= sub_wire22(28);
	sub_wire1(42, 29)    <= sub_wire22(29);
	sub_wire1(42, 30)    <= sub_wire22(30);
	sub_wire1(42, 31)    <= sub_wire22(31);
	sub_wire1(41, 0)    <= sub_wire23(0);
	sub_wire1(41, 1)    <= sub_wire23(1);
	sub_wire1(41, 2)    <= sub_wire23(2);
	sub_wire1(41, 3)    <= sub_wire23(3);
	sub_wire1(41, 4)    <= sub_wire23(4);
	sub_wire1(41, 5)    <= sub_wire23(5);
	sub_wire1(41, 6)    <= sub_wire23(6);
	sub_wire1(41, 7)    <= sub_wire23(7);
	sub_wire1(41, 8)    <= sub_wire23(8);
	sub_wire1(41, 9)    <= sub_wire23(9);
	sub_wire1(41, 10)    <= sub_wire23(10);
	sub_wire1(41, 11)    <= sub_wire23(11);
	sub_wire1(41, 12)    <= sub_wire23(12);
	sub_wire1(41, 13)    <= sub_wire23(13);
	sub_wire1(41, 14)    <= sub_wire23(14);
	sub_wire1(41, 15)    <= sub_wire23(15);
	sub_wire1(41, 16)    <= sub_wire23(16);
	sub_wire1(41, 17)    <= sub_wire23(17);
	sub_wire1(41, 18)    <= sub_wire23(18);
	sub_wire1(41, 19)    <= sub_wire23(19);
	sub_wire1(41, 20)    <= sub_wire23(20);
	sub_wire1(41, 21)    <= sub_wire23(21);
	sub_wire1(41, 22)    <= sub_wire23(22);
	sub_wire1(41, 23)    <= sub_wire23(23);
	sub_wire1(41, 24)    <= sub_wire23(24);
	sub_wire1(41, 25)    <= sub_wire23(25);
	sub_wire1(41, 26)    <= sub_wire23(26);
	sub_wire1(41, 27)    <= sub_wire23(27);
	sub_wire1(41, 28)    <= sub_wire23(28);
	sub_wire1(41, 29)    <= sub_wire23(29);
	sub_wire1(41, 30)    <= sub_wire23(30);
	sub_wire1(41, 31)    <= sub_wire23(31);
	sub_wire1(40, 0)    <= sub_wire24(0);
	sub_wire1(40, 1)    <= sub_wire24(1);
	sub_wire1(40, 2)    <= sub_wire24(2);
	sub_wire1(40, 3)    <= sub_wire24(3);
	sub_wire1(40, 4)    <= sub_wire24(4);
	sub_wire1(40, 5)    <= sub_wire24(5);
	sub_wire1(40, 6)    <= sub_wire24(6);
	sub_wire1(40, 7)    <= sub_wire24(7);
	sub_wire1(40, 8)    <= sub_wire24(8);
	sub_wire1(40, 9)    <= sub_wire24(9);
	sub_wire1(40, 10)    <= sub_wire24(10);
	sub_wire1(40, 11)    <= sub_wire24(11);
	sub_wire1(40, 12)    <= sub_wire24(12);
	sub_wire1(40, 13)    <= sub_wire24(13);
	sub_wire1(40, 14)    <= sub_wire24(14);
	sub_wire1(40, 15)    <= sub_wire24(15);
	sub_wire1(40, 16)    <= sub_wire24(16);
	sub_wire1(40, 17)    <= sub_wire24(17);
	sub_wire1(40, 18)    <= sub_wire24(18);
	sub_wire1(40, 19)    <= sub_wire24(19);
	sub_wire1(40, 20)    <= sub_wire24(20);
	sub_wire1(40, 21)    <= sub_wire24(21);
	sub_wire1(40, 22)    <= sub_wire24(22);
	sub_wire1(40, 23)    <= sub_wire24(23);
	sub_wire1(40, 24)    <= sub_wire24(24);
	sub_wire1(40, 25)    <= sub_wire24(25);
	sub_wire1(40, 26)    <= sub_wire24(26);
	sub_wire1(40, 27)    <= sub_wire24(27);
	sub_wire1(40, 28)    <= sub_wire24(28);
	sub_wire1(40, 29)    <= sub_wire24(29);
	sub_wire1(40, 30)    <= sub_wire24(30);
	sub_wire1(40, 31)    <= sub_wire24(31);
	sub_wire1(39, 0)    <= sub_wire25(0);
	sub_wire1(39, 1)    <= sub_wire25(1);
	sub_wire1(39, 2)    <= sub_wire25(2);
	sub_wire1(39, 3)    <= sub_wire25(3);
	sub_wire1(39, 4)    <= sub_wire25(4);
	sub_wire1(39, 5)    <= sub_wire25(5);
	sub_wire1(39, 6)    <= sub_wire25(6);
	sub_wire1(39, 7)    <= sub_wire25(7);
	sub_wire1(39, 8)    <= sub_wire25(8);
	sub_wire1(39, 9)    <= sub_wire25(9);
	sub_wire1(39, 10)    <= sub_wire25(10);
	sub_wire1(39, 11)    <= sub_wire25(11);
	sub_wire1(39, 12)    <= sub_wire25(12);
	sub_wire1(39, 13)    <= sub_wire25(13);
	sub_wire1(39, 14)    <= sub_wire25(14);
	sub_wire1(39, 15)    <= sub_wire25(15);
	sub_wire1(39, 16)    <= sub_wire25(16);
	sub_wire1(39, 17)    <= sub_wire25(17);
	sub_wire1(39, 18)    <= sub_wire25(18);
	sub_wire1(39, 19)    <= sub_wire25(19);
	sub_wire1(39, 20)    <= sub_wire25(20);
	sub_wire1(39, 21)    <= sub_wire25(21);
	sub_wire1(39, 22)    <= sub_wire25(22);
	sub_wire1(39, 23)    <= sub_wire25(23);
	sub_wire1(39, 24)    <= sub_wire25(24);
	sub_wire1(39, 25)    <= sub_wire25(25);
	sub_wire1(39, 26)    <= sub_wire25(26);
	sub_wire1(39, 27)    <= sub_wire25(27);
	sub_wire1(39, 28)    <= sub_wire25(28);
	sub_wire1(39, 29)    <= sub_wire25(29);
	sub_wire1(39, 30)    <= sub_wire25(30);
	sub_wire1(39, 31)    <= sub_wire25(31);
	sub_wire1(38, 0)    <= sub_wire26(0);
	sub_wire1(38, 1)    <= sub_wire26(1);
	sub_wire1(38, 2)    <= sub_wire26(2);
	sub_wire1(38, 3)    <= sub_wire26(3);
	sub_wire1(38, 4)    <= sub_wire26(4);
	sub_wire1(38, 5)    <= sub_wire26(5);
	sub_wire1(38, 6)    <= sub_wire26(6);
	sub_wire1(38, 7)    <= sub_wire26(7);
	sub_wire1(38, 8)    <= sub_wire26(8);
	sub_wire1(38, 9)    <= sub_wire26(9);
	sub_wire1(38, 10)    <= sub_wire26(10);
	sub_wire1(38, 11)    <= sub_wire26(11);
	sub_wire1(38, 12)    <= sub_wire26(12);
	sub_wire1(38, 13)    <= sub_wire26(13);
	sub_wire1(38, 14)    <= sub_wire26(14);
	sub_wire1(38, 15)    <= sub_wire26(15);
	sub_wire1(38, 16)    <= sub_wire26(16);
	sub_wire1(38, 17)    <= sub_wire26(17);
	sub_wire1(38, 18)    <= sub_wire26(18);
	sub_wire1(38, 19)    <= sub_wire26(19);
	sub_wire1(38, 20)    <= sub_wire26(20);
	sub_wire1(38, 21)    <= sub_wire26(21);
	sub_wire1(38, 22)    <= sub_wire26(22);
	sub_wire1(38, 23)    <= sub_wire26(23);
	sub_wire1(38, 24)    <= sub_wire26(24);
	sub_wire1(38, 25)    <= sub_wire26(25);
	sub_wire1(38, 26)    <= sub_wire26(26);
	sub_wire1(38, 27)    <= sub_wire26(27);
	sub_wire1(38, 28)    <= sub_wire26(28);
	sub_wire1(38, 29)    <= sub_wire26(29);
	sub_wire1(38, 30)    <= sub_wire26(30);
	sub_wire1(38, 31)    <= sub_wire26(31);
	sub_wire1(37, 0)    <= sub_wire27(0);
	sub_wire1(37, 1)    <= sub_wire27(1);
	sub_wire1(37, 2)    <= sub_wire27(2);
	sub_wire1(37, 3)    <= sub_wire27(3);
	sub_wire1(37, 4)    <= sub_wire27(4);
	sub_wire1(37, 5)    <= sub_wire27(5);
	sub_wire1(37, 6)    <= sub_wire27(6);
	sub_wire1(37, 7)    <= sub_wire27(7);
	sub_wire1(37, 8)    <= sub_wire27(8);
	sub_wire1(37, 9)    <= sub_wire27(9);
	sub_wire1(37, 10)    <= sub_wire27(10);
	sub_wire1(37, 11)    <= sub_wire27(11);
	sub_wire1(37, 12)    <= sub_wire27(12);
	sub_wire1(37, 13)    <= sub_wire27(13);
	sub_wire1(37, 14)    <= sub_wire27(14);
	sub_wire1(37, 15)    <= sub_wire27(15);
	sub_wire1(37, 16)    <= sub_wire27(16);
	sub_wire1(37, 17)    <= sub_wire27(17);
	sub_wire1(37, 18)    <= sub_wire27(18);
	sub_wire1(37, 19)    <= sub_wire27(19);
	sub_wire1(37, 20)    <= sub_wire27(20);
	sub_wire1(37, 21)    <= sub_wire27(21);
	sub_wire1(37, 22)    <= sub_wire27(22);
	sub_wire1(37, 23)    <= sub_wire27(23);
	sub_wire1(37, 24)    <= sub_wire27(24);
	sub_wire1(37, 25)    <= sub_wire27(25);
	sub_wire1(37, 26)    <= sub_wire27(26);
	sub_wire1(37, 27)    <= sub_wire27(27);
	sub_wire1(37, 28)    <= sub_wire27(28);
	sub_wire1(37, 29)    <= sub_wire27(29);
	sub_wire1(37, 30)    <= sub_wire27(30);
	sub_wire1(37, 31)    <= sub_wire27(31);
	sub_wire1(36, 0)    <= sub_wire28(0);
	sub_wire1(36, 1)    <= sub_wire28(1);
	sub_wire1(36, 2)    <= sub_wire28(2);
	sub_wire1(36, 3)    <= sub_wire28(3);
	sub_wire1(36, 4)    <= sub_wire28(4);
	sub_wire1(36, 5)    <= sub_wire28(5);
	sub_wire1(36, 6)    <= sub_wire28(6);
	sub_wire1(36, 7)    <= sub_wire28(7);
	sub_wire1(36, 8)    <= sub_wire28(8);
	sub_wire1(36, 9)    <= sub_wire28(9);
	sub_wire1(36, 10)    <= sub_wire28(10);
	sub_wire1(36, 11)    <= sub_wire28(11);
	sub_wire1(36, 12)    <= sub_wire28(12);
	sub_wire1(36, 13)    <= sub_wire28(13);
	sub_wire1(36, 14)    <= sub_wire28(14);
	sub_wire1(36, 15)    <= sub_wire28(15);
	sub_wire1(36, 16)    <= sub_wire28(16);
	sub_wire1(36, 17)    <= sub_wire28(17);
	sub_wire1(36, 18)    <= sub_wire28(18);
	sub_wire1(36, 19)    <= sub_wire28(19);
	sub_wire1(36, 20)    <= sub_wire28(20);
	sub_wire1(36, 21)    <= sub_wire28(21);
	sub_wire1(36, 22)    <= sub_wire28(22);
	sub_wire1(36, 23)    <= sub_wire28(23);
	sub_wire1(36, 24)    <= sub_wire28(24);
	sub_wire1(36, 25)    <= sub_wire28(25);
	sub_wire1(36, 26)    <= sub_wire28(26);
	sub_wire1(36, 27)    <= sub_wire28(27);
	sub_wire1(36, 28)    <= sub_wire28(28);
	sub_wire1(36, 29)    <= sub_wire28(29);
	sub_wire1(36, 30)    <= sub_wire28(30);
	sub_wire1(36, 31)    <= sub_wire28(31);
	sub_wire1(35, 0)    <= sub_wire29(0);
	sub_wire1(35, 1)    <= sub_wire29(1);
	sub_wire1(35, 2)    <= sub_wire29(2);
	sub_wire1(35, 3)    <= sub_wire29(3);
	sub_wire1(35, 4)    <= sub_wire29(4);
	sub_wire1(35, 5)    <= sub_wire29(5);
	sub_wire1(35, 6)    <= sub_wire29(6);
	sub_wire1(35, 7)    <= sub_wire29(7);
	sub_wire1(35, 8)    <= sub_wire29(8);
	sub_wire1(35, 9)    <= sub_wire29(9);
	sub_wire1(35, 10)    <= sub_wire29(10);
	sub_wire1(35, 11)    <= sub_wire29(11);
	sub_wire1(35, 12)    <= sub_wire29(12);
	sub_wire1(35, 13)    <= sub_wire29(13);
	sub_wire1(35, 14)    <= sub_wire29(14);
	sub_wire1(35, 15)    <= sub_wire29(15);
	sub_wire1(35, 16)    <= sub_wire29(16);
	sub_wire1(35, 17)    <= sub_wire29(17);
	sub_wire1(35, 18)    <= sub_wire29(18);
	sub_wire1(35, 19)    <= sub_wire29(19);
	sub_wire1(35, 20)    <= sub_wire29(20);
	sub_wire1(35, 21)    <= sub_wire29(21);
	sub_wire1(35, 22)    <= sub_wire29(22);
	sub_wire1(35, 23)    <= sub_wire29(23);
	sub_wire1(35, 24)    <= sub_wire29(24);
	sub_wire1(35, 25)    <= sub_wire29(25);
	sub_wire1(35, 26)    <= sub_wire29(26);
	sub_wire1(35, 27)    <= sub_wire29(27);
	sub_wire1(35, 28)    <= sub_wire29(28);
	sub_wire1(35, 29)    <= sub_wire29(29);
	sub_wire1(35, 30)    <= sub_wire29(30);
	sub_wire1(35, 31)    <= sub_wire29(31);
	sub_wire1(34, 0)    <= sub_wire30(0);
	sub_wire1(34, 1)    <= sub_wire30(1);
	sub_wire1(34, 2)    <= sub_wire30(2);
	sub_wire1(34, 3)    <= sub_wire30(3);
	sub_wire1(34, 4)    <= sub_wire30(4);
	sub_wire1(34, 5)    <= sub_wire30(5);
	sub_wire1(34, 6)    <= sub_wire30(6);
	sub_wire1(34, 7)    <= sub_wire30(7);
	sub_wire1(34, 8)    <= sub_wire30(8);
	sub_wire1(34, 9)    <= sub_wire30(9);
	sub_wire1(34, 10)    <= sub_wire30(10);
	sub_wire1(34, 11)    <= sub_wire30(11);
	sub_wire1(34, 12)    <= sub_wire30(12);
	sub_wire1(34, 13)    <= sub_wire30(13);
	sub_wire1(34, 14)    <= sub_wire30(14);
	sub_wire1(34, 15)    <= sub_wire30(15);
	sub_wire1(34, 16)    <= sub_wire30(16);
	sub_wire1(34, 17)    <= sub_wire30(17);
	sub_wire1(34, 18)    <= sub_wire30(18);
	sub_wire1(34, 19)    <= sub_wire30(19);
	sub_wire1(34, 20)    <= sub_wire30(20);
	sub_wire1(34, 21)    <= sub_wire30(21);
	sub_wire1(34, 22)    <= sub_wire30(22);
	sub_wire1(34, 23)    <= sub_wire30(23);
	sub_wire1(34, 24)    <= sub_wire30(24);
	sub_wire1(34, 25)    <= sub_wire30(25);
	sub_wire1(34, 26)    <= sub_wire30(26);
	sub_wire1(34, 27)    <= sub_wire30(27);
	sub_wire1(34, 28)    <= sub_wire30(28);
	sub_wire1(34, 29)    <= sub_wire30(29);
	sub_wire1(34, 30)    <= sub_wire30(30);
	sub_wire1(34, 31)    <= sub_wire30(31);
	sub_wire1(33, 0)    <= sub_wire31(0);
	sub_wire1(33, 1)    <= sub_wire31(1);
	sub_wire1(33, 2)    <= sub_wire31(2);
	sub_wire1(33, 3)    <= sub_wire31(3);
	sub_wire1(33, 4)    <= sub_wire31(4);
	sub_wire1(33, 5)    <= sub_wire31(5);
	sub_wire1(33, 6)    <= sub_wire31(6);
	sub_wire1(33, 7)    <= sub_wire31(7);
	sub_wire1(33, 8)    <= sub_wire31(8);
	sub_wire1(33, 9)    <= sub_wire31(9);
	sub_wire1(33, 10)    <= sub_wire31(10);
	sub_wire1(33, 11)    <= sub_wire31(11);
	sub_wire1(33, 12)    <= sub_wire31(12);
	sub_wire1(33, 13)    <= sub_wire31(13);
	sub_wire1(33, 14)    <= sub_wire31(14);
	sub_wire1(33, 15)    <= sub_wire31(15);
	sub_wire1(33, 16)    <= sub_wire31(16);
	sub_wire1(33, 17)    <= sub_wire31(17);
	sub_wire1(33, 18)    <= sub_wire31(18);
	sub_wire1(33, 19)    <= sub_wire31(19);
	sub_wire1(33, 20)    <= sub_wire31(20);
	sub_wire1(33, 21)    <= sub_wire31(21);
	sub_wire1(33, 22)    <= sub_wire31(22);
	sub_wire1(33, 23)    <= sub_wire31(23);
	sub_wire1(33, 24)    <= sub_wire31(24);
	sub_wire1(33, 25)    <= sub_wire31(25);
	sub_wire1(33, 26)    <= sub_wire31(26);
	sub_wire1(33, 27)    <= sub_wire31(27);
	sub_wire1(33, 28)    <= sub_wire31(28);
	sub_wire1(33, 29)    <= sub_wire31(29);
	sub_wire1(33, 30)    <= sub_wire31(30);
	sub_wire1(33, 31)    <= sub_wire31(31);
	sub_wire1(32, 0)    <= sub_wire32(0);
	sub_wire1(32, 1)    <= sub_wire32(1);
	sub_wire1(32, 2)    <= sub_wire32(2);
	sub_wire1(32, 3)    <= sub_wire32(3);
	sub_wire1(32, 4)    <= sub_wire32(4);
	sub_wire1(32, 5)    <= sub_wire32(5);
	sub_wire1(32, 6)    <= sub_wire32(6);
	sub_wire1(32, 7)    <= sub_wire32(7);
	sub_wire1(32, 8)    <= sub_wire32(8);
	sub_wire1(32, 9)    <= sub_wire32(9);
	sub_wire1(32, 10)    <= sub_wire32(10);
	sub_wire1(32, 11)    <= sub_wire32(11);
	sub_wire1(32, 12)    <= sub_wire32(12);
	sub_wire1(32, 13)    <= sub_wire32(13);
	sub_wire1(32, 14)    <= sub_wire32(14);
	sub_wire1(32, 15)    <= sub_wire32(15);
	sub_wire1(32, 16)    <= sub_wire32(16);
	sub_wire1(32, 17)    <= sub_wire32(17);
	sub_wire1(32, 18)    <= sub_wire32(18);
	sub_wire1(32, 19)    <= sub_wire32(19);
	sub_wire1(32, 20)    <= sub_wire32(20);
	sub_wire1(32, 21)    <= sub_wire32(21);
	sub_wire1(32, 22)    <= sub_wire32(22);
	sub_wire1(32, 23)    <= sub_wire32(23);
	sub_wire1(32, 24)    <= sub_wire32(24);
	sub_wire1(32, 25)    <= sub_wire32(25);
	sub_wire1(32, 26)    <= sub_wire32(26);
	sub_wire1(32, 27)    <= sub_wire32(27);
	sub_wire1(32, 28)    <= sub_wire32(28);
	sub_wire1(32, 29)    <= sub_wire32(29);
	sub_wire1(32, 30)    <= sub_wire32(30);
	sub_wire1(32, 31)    <= sub_wire32(31);
	sub_wire1(31, 0)    <= sub_wire33(0);
	sub_wire1(31, 1)    <= sub_wire33(1);
	sub_wire1(31, 2)    <= sub_wire33(2);
	sub_wire1(31, 3)    <= sub_wire33(3);
	sub_wire1(31, 4)    <= sub_wire33(4);
	sub_wire1(31, 5)    <= sub_wire33(5);
	sub_wire1(31, 6)    <= sub_wire33(6);
	sub_wire1(31, 7)    <= sub_wire33(7);
	sub_wire1(31, 8)    <= sub_wire33(8);
	sub_wire1(31, 9)    <= sub_wire33(9);
	sub_wire1(31, 10)    <= sub_wire33(10);
	sub_wire1(31, 11)    <= sub_wire33(11);
	sub_wire1(31, 12)    <= sub_wire33(12);
	sub_wire1(31, 13)    <= sub_wire33(13);
	sub_wire1(31, 14)    <= sub_wire33(14);
	sub_wire1(31, 15)    <= sub_wire33(15);
	sub_wire1(31, 16)    <= sub_wire33(16);
	sub_wire1(31, 17)    <= sub_wire33(17);
	sub_wire1(31, 18)    <= sub_wire33(18);
	sub_wire1(31, 19)    <= sub_wire33(19);
	sub_wire1(31, 20)    <= sub_wire33(20);
	sub_wire1(31, 21)    <= sub_wire33(21);
	sub_wire1(31, 22)    <= sub_wire33(22);
	sub_wire1(31, 23)    <= sub_wire33(23);
	sub_wire1(31, 24)    <= sub_wire33(24);
	sub_wire1(31, 25)    <= sub_wire33(25);
	sub_wire1(31, 26)    <= sub_wire33(26);
	sub_wire1(31, 27)    <= sub_wire33(27);
	sub_wire1(31, 28)    <= sub_wire33(28);
	sub_wire1(31, 29)    <= sub_wire33(29);
	sub_wire1(31, 30)    <= sub_wire33(30);
	sub_wire1(31, 31)    <= sub_wire33(31);
	sub_wire1(30, 0)    <= sub_wire34(0);
	sub_wire1(30, 1)    <= sub_wire34(1);
	sub_wire1(30, 2)    <= sub_wire34(2);
	sub_wire1(30, 3)    <= sub_wire34(3);
	sub_wire1(30, 4)    <= sub_wire34(4);
	sub_wire1(30, 5)    <= sub_wire34(5);
	sub_wire1(30, 6)    <= sub_wire34(6);
	sub_wire1(30, 7)    <= sub_wire34(7);
	sub_wire1(30, 8)    <= sub_wire34(8);
	sub_wire1(30, 9)    <= sub_wire34(9);
	sub_wire1(30, 10)    <= sub_wire34(10);
	sub_wire1(30, 11)    <= sub_wire34(11);
	sub_wire1(30, 12)    <= sub_wire34(12);
	sub_wire1(30, 13)    <= sub_wire34(13);
	sub_wire1(30, 14)    <= sub_wire34(14);
	sub_wire1(30, 15)    <= sub_wire34(15);
	sub_wire1(30, 16)    <= sub_wire34(16);
	sub_wire1(30, 17)    <= sub_wire34(17);
	sub_wire1(30, 18)    <= sub_wire34(18);
	sub_wire1(30, 19)    <= sub_wire34(19);
	sub_wire1(30, 20)    <= sub_wire34(20);
	sub_wire1(30, 21)    <= sub_wire34(21);
	sub_wire1(30, 22)    <= sub_wire34(22);
	sub_wire1(30, 23)    <= sub_wire34(23);
	sub_wire1(30, 24)    <= sub_wire34(24);
	sub_wire1(30, 25)    <= sub_wire34(25);
	sub_wire1(30, 26)    <= sub_wire34(26);
	sub_wire1(30, 27)    <= sub_wire34(27);
	sub_wire1(30, 28)    <= sub_wire34(28);
	sub_wire1(30, 29)    <= sub_wire34(29);
	sub_wire1(30, 30)    <= sub_wire34(30);
	sub_wire1(30, 31)    <= sub_wire34(31);
	sub_wire1(29, 0)    <= sub_wire35(0);
	sub_wire1(29, 1)    <= sub_wire35(1);
	sub_wire1(29, 2)    <= sub_wire35(2);
	sub_wire1(29, 3)    <= sub_wire35(3);
	sub_wire1(29, 4)    <= sub_wire35(4);
	sub_wire1(29, 5)    <= sub_wire35(5);
	sub_wire1(29, 6)    <= sub_wire35(6);
	sub_wire1(29, 7)    <= sub_wire35(7);
	sub_wire1(29, 8)    <= sub_wire35(8);
	sub_wire1(29, 9)    <= sub_wire35(9);
	sub_wire1(29, 10)    <= sub_wire35(10);
	sub_wire1(29, 11)    <= sub_wire35(11);
	sub_wire1(29, 12)    <= sub_wire35(12);
	sub_wire1(29, 13)    <= sub_wire35(13);
	sub_wire1(29, 14)    <= sub_wire35(14);
	sub_wire1(29, 15)    <= sub_wire35(15);
	sub_wire1(29, 16)    <= sub_wire35(16);
	sub_wire1(29, 17)    <= sub_wire35(17);
	sub_wire1(29, 18)    <= sub_wire35(18);
	sub_wire1(29, 19)    <= sub_wire35(19);
	sub_wire1(29, 20)    <= sub_wire35(20);
	sub_wire1(29, 21)    <= sub_wire35(21);
	sub_wire1(29, 22)    <= sub_wire35(22);
	sub_wire1(29, 23)    <= sub_wire35(23);
	sub_wire1(29, 24)    <= sub_wire35(24);
	sub_wire1(29, 25)    <= sub_wire35(25);
	sub_wire1(29, 26)    <= sub_wire35(26);
	sub_wire1(29, 27)    <= sub_wire35(27);
	sub_wire1(29, 28)    <= sub_wire35(28);
	sub_wire1(29, 29)    <= sub_wire35(29);
	sub_wire1(29, 30)    <= sub_wire35(30);
	sub_wire1(29, 31)    <= sub_wire35(31);
	sub_wire1(28, 0)    <= sub_wire36(0);
	sub_wire1(28, 1)    <= sub_wire36(1);
	sub_wire1(28, 2)    <= sub_wire36(2);
	sub_wire1(28, 3)    <= sub_wire36(3);
	sub_wire1(28, 4)    <= sub_wire36(4);
	sub_wire1(28, 5)    <= sub_wire36(5);
	sub_wire1(28, 6)    <= sub_wire36(6);
	sub_wire1(28, 7)    <= sub_wire36(7);
	sub_wire1(28, 8)    <= sub_wire36(8);
	sub_wire1(28, 9)    <= sub_wire36(9);
	sub_wire1(28, 10)    <= sub_wire36(10);
	sub_wire1(28, 11)    <= sub_wire36(11);
	sub_wire1(28, 12)    <= sub_wire36(12);
	sub_wire1(28, 13)    <= sub_wire36(13);
	sub_wire1(28, 14)    <= sub_wire36(14);
	sub_wire1(28, 15)    <= sub_wire36(15);
	sub_wire1(28, 16)    <= sub_wire36(16);
	sub_wire1(28, 17)    <= sub_wire36(17);
	sub_wire1(28, 18)    <= sub_wire36(18);
	sub_wire1(28, 19)    <= sub_wire36(19);
	sub_wire1(28, 20)    <= sub_wire36(20);
	sub_wire1(28, 21)    <= sub_wire36(21);
	sub_wire1(28, 22)    <= sub_wire36(22);
	sub_wire1(28, 23)    <= sub_wire36(23);
	sub_wire1(28, 24)    <= sub_wire36(24);
	sub_wire1(28, 25)    <= sub_wire36(25);
	sub_wire1(28, 26)    <= sub_wire36(26);
	sub_wire1(28, 27)    <= sub_wire36(27);
	sub_wire1(28, 28)    <= sub_wire36(28);
	sub_wire1(28, 29)    <= sub_wire36(29);
	sub_wire1(28, 30)    <= sub_wire36(30);
	sub_wire1(28, 31)    <= sub_wire36(31);
	sub_wire1(27, 0)    <= sub_wire37(0);
	sub_wire1(27, 1)    <= sub_wire37(1);
	sub_wire1(27, 2)    <= sub_wire37(2);
	sub_wire1(27, 3)    <= sub_wire37(3);
	sub_wire1(27, 4)    <= sub_wire37(4);
	sub_wire1(27, 5)    <= sub_wire37(5);
	sub_wire1(27, 6)    <= sub_wire37(6);
	sub_wire1(27, 7)    <= sub_wire37(7);
	sub_wire1(27, 8)    <= sub_wire37(8);
	sub_wire1(27, 9)    <= sub_wire37(9);
	sub_wire1(27, 10)    <= sub_wire37(10);
	sub_wire1(27, 11)    <= sub_wire37(11);
	sub_wire1(27, 12)    <= sub_wire37(12);
	sub_wire1(27, 13)    <= sub_wire37(13);
	sub_wire1(27, 14)    <= sub_wire37(14);
	sub_wire1(27, 15)    <= sub_wire37(15);
	sub_wire1(27, 16)    <= sub_wire37(16);
	sub_wire1(27, 17)    <= sub_wire37(17);
	sub_wire1(27, 18)    <= sub_wire37(18);
	sub_wire1(27, 19)    <= sub_wire37(19);
	sub_wire1(27, 20)    <= sub_wire37(20);
	sub_wire1(27, 21)    <= sub_wire37(21);
	sub_wire1(27, 22)    <= sub_wire37(22);
	sub_wire1(27, 23)    <= sub_wire37(23);
	sub_wire1(27, 24)    <= sub_wire37(24);
	sub_wire1(27, 25)    <= sub_wire37(25);
	sub_wire1(27, 26)    <= sub_wire37(26);
	sub_wire1(27, 27)    <= sub_wire37(27);
	sub_wire1(27, 28)    <= sub_wire37(28);
	sub_wire1(27, 29)    <= sub_wire37(29);
	sub_wire1(27, 30)    <= sub_wire37(30);
	sub_wire1(27, 31)    <= sub_wire37(31);
	sub_wire1(26, 0)    <= sub_wire38(0);
	sub_wire1(26, 1)    <= sub_wire38(1);
	sub_wire1(26, 2)    <= sub_wire38(2);
	sub_wire1(26, 3)    <= sub_wire38(3);
	sub_wire1(26, 4)    <= sub_wire38(4);
	sub_wire1(26, 5)    <= sub_wire38(5);
	sub_wire1(26, 6)    <= sub_wire38(6);
	sub_wire1(26, 7)    <= sub_wire38(7);
	sub_wire1(26, 8)    <= sub_wire38(8);
	sub_wire1(26, 9)    <= sub_wire38(9);
	sub_wire1(26, 10)    <= sub_wire38(10);
	sub_wire1(26, 11)    <= sub_wire38(11);
	sub_wire1(26, 12)    <= sub_wire38(12);
	sub_wire1(26, 13)    <= sub_wire38(13);
	sub_wire1(26, 14)    <= sub_wire38(14);
	sub_wire1(26, 15)    <= sub_wire38(15);
	sub_wire1(26, 16)    <= sub_wire38(16);
	sub_wire1(26, 17)    <= sub_wire38(17);
	sub_wire1(26, 18)    <= sub_wire38(18);
	sub_wire1(26, 19)    <= sub_wire38(19);
	sub_wire1(26, 20)    <= sub_wire38(20);
	sub_wire1(26, 21)    <= sub_wire38(21);
	sub_wire1(26, 22)    <= sub_wire38(22);
	sub_wire1(26, 23)    <= sub_wire38(23);
	sub_wire1(26, 24)    <= sub_wire38(24);
	sub_wire1(26, 25)    <= sub_wire38(25);
	sub_wire1(26, 26)    <= sub_wire38(26);
	sub_wire1(26, 27)    <= sub_wire38(27);
	sub_wire1(26, 28)    <= sub_wire38(28);
	sub_wire1(26, 29)    <= sub_wire38(29);
	sub_wire1(26, 30)    <= sub_wire38(30);
	sub_wire1(26, 31)    <= sub_wire38(31);
	sub_wire1(25, 0)    <= sub_wire39(0);
	sub_wire1(25, 1)    <= sub_wire39(1);
	sub_wire1(25, 2)    <= sub_wire39(2);
	sub_wire1(25, 3)    <= sub_wire39(3);
	sub_wire1(25, 4)    <= sub_wire39(4);
	sub_wire1(25, 5)    <= sub_wire39(5);
	sub_wire1(25, 6)    <= sub_wire39(6);
	sub_wire1(25, 7)    <= sub_wire39(7);
	sub_wire1(25, 8)    <= sub_wire39(8);
	sub_wire1(25, 9)    <= sub_wire39(9);
	sub_wire1(25, 10)    <= sub_wire39(10);
	sub_wire1(25, 11)    <= sub_wire39(11);
	sub_wire1(25, 12)    <= sub_wire39(12);
	sub_wire1(25, 13)    <= sub_wire39(13);
	sub_wire1(25, 14)    <= sub_wire39(14);
	sub_wire1(25, 15)    <= sub_wire39(15);
	sub_wire1(25, 16)    <= sub_wire39(16);
	sub_wire1(25, 17)    <= sub_wire39(17);
	sub_wire1(25, 18)    <= sub_wire39(18);
	sub_wire1(25, 19)    <= sub_wire39(19);
	sub_wire1(25, 20)    <= sub_wire39(20);
	sub_wire1(25, 21)    <= sub_wire39(21);
	sub_wire1(25, 22)    <= sub_wire39(22);
	sub_wire1(25, 23)    <= sub_wire39(23);
	sub_wire1(25, 24)    <= sub_wire39(24);
	sub_wire1(25, 25)    <= sub_wire39(25);
	sub_wire1(25, 26)    <= sub_wire39(26);
	sub_wire1(25, 27)    <= sub_wire39(27);
	sub_wire1(25, 28)    <= sub_wire39(28);
	sub_wire1(25, 29)    <= sub_wire39(29);
	sub_wire1(25, 30)    <= sub_wire39(30);
	sub_wire1(25, 31)    <= sub_wire39(31);
	sub_wire1(24, 0)    <= sub_wire40(0);
	sub_wire1(24, 1)    <= sub_wire40(1);
	sub_wire1(24, 2)    <= sub_wire40(2);
	sub_wire1(24, 3)    <= sub_wire40(3);
	sub_wire1(24, 4)    <= sub_wire40(4);
	sub_wire1(24, 5)    <= sub_wire40(5);
	sub_wire1(24, 6)    <= sub_wire40(6);
	sub_wire1(24, 7)    <= sub_wire40(7);
	sub_wire1(24, 8)    <= sub_wire40(8);
	sub_wire1(24, 9)    <= sub_wire40(9);
	sub_wire1(24, 10)    <= sub_wire40(10);
	sub_wire1(24, 11)    <= sub_wire40(11);
	sub_wire1(24, 12)    <= sub_wire40(12);
	sub_wire1(24, 13)    <= sub_wire40(13);
	sub_wire1(24, 14)    <= sub_wire40(14);
	sub_wire1(24, 15)    <= sub_wire40(15);
	sub_wire1(24, 16)    <= sub_wire40(16);
	sub_wire1(24, 17)    <= sub_wire40(17);
	sub_wire1(24, 18)    <= sub_wire40(18);
	sub_wire1(24, 19)    <= sub_wire40(19);
	sub_wire1(24, 20)    <= sub_wire40(20);
	sub_wire1(24, 21)    <= sub_wire40(21);
	sub_wire1(24, 22)    <= sub_wire40(22);
	sub_wire1(24, 23)    <= sub_wire40(23);
	sub_wire1(24, 24)    <= sub_wire40(24);
	sub_wire1(24, 25)    <= sub_wire40(25);
	sub_wire1(24, 26)    <= sub_wire40(26);
	sub_wire1(24, 27)    <= sub_wire40(27);
	sub_wire1(24, 28)    <= sub_wire40(28);
	sub_wire1(24, 29)    <= sub_wire40(29);
	sub_wire1(24, 30)    <= sub_wire40(30);
	sub_wire1(24, 31)    <= sub_wire40(31);
	sub_wire1(23, 0)    <= sub_wire41(0);
	sub_wire1(23, 1)    <= sub_wire41(1);
	sub_wire1(23, 2)    <= sub_wire41(2);
	sub_wire1(23, 3)    <= sub_wire41(3);
	sub_wire1(23, 4)    <= sub_wire41(4);
	sub_wire1(23, 5)    <= sub_wire41(5);
	sub_wire1(23, 6)    <= sub_wire41(6);
	sub_wire1(23, 7)    <= sub_wire41(7);
	sub_wire1(23, 8)    <= sub_wire41(8);
	sub_wire1(23, 9)    <= sub_wire41(9);
	sub_wire1(23, 10)    <= sub_wire41(10);
	sub_wire1(23, 11)    <= sub_wire41(11);
	sub_wire1(23, 12)    <= sub_wire41(12);
	sub_wire1(23, 13)    <= sub_wire41(13);
	sub_wire1(23, 14)    <= sub_wire41(14);
	sub_wire1(23, 15)    <= sub_wire41(15);
	sub_wire1(23, 16)    <= sub_wire41(16);
	sub_wire1(23, 17)    <= sub_wire41(17);
	sub_wire1(23, 18)    <= sub_wire41(18);
	sub_wire1(23, 19)    <= sub_wire41(19);
	sub_wire1(23, 20)    <= sub_wire41(20);
	sub_wire1(23, 21)    <= sub_wire41(21);
	sub_wire1(23, 22)    <= sub_wire41(22);
	sub_wire1(23, 23)    <= sub_wire41(23);
	sub_wire1(23, 24)    <= sub_wire41(24);
	sub_wire1(23, 25)    <= sub_wire41(25);
	sub_wire1(23, 26)    <= sub_wire41(26);
	sub_wire1(23, 27)    <= sub_wire41(27);
	sub_wire1(23, 28)    <= sub_wire41(28);
	sub_wire1(23, 29)    <= sub_wire41(29);
	sub_wire1(23, 30)    <= sub_wire41(30);
	sub_wire1(23, 31)    <= sub_wire41(31);
	sub_wire1(22, 0)    <= sub_wire42(0);
	sub_wire1(22, 1)    <= sub_wire42(1);
	sub_wire1(22, 2)    <= sub_wire42(2);
	sub_wire1(22, 3)    <= sub_wire42(3);
	sub_wire1(22, 4)    <= sub_wire42(4);
	sub_wire1(22, 5)    <= sub_wire42(5);
	sub_wire1(22, 6)    <= sub_wire42(6);
	sub_wire1(22, 7)    <= sub_wire42(7);
	sub_wire1(22, 8)    <= sub_wire42(8);
	sub_wire1(22, 9)    <= sub_wire42(9);
	sub_wire1(22, 10)    <= sub_wire42(10);
	sub_wire1(22, 11)    <= sub_wire42(11);
	sub_wire1(22, 12)    <= sub_wire42(12);
	sub_wire1(22, 13)    <= sub_wire42(13);
	sub_wire1(22, 14)    <= sub_wire42(14);
	sub_wire1(22, 15)    <= sub_wire42(15);
	sub_wire1(22, 16)    <= sub_wire42(16);
	sub_wire1(22, 17)    <= sub_wire42(17);
	sub_wire1(22, 18)    <= sub_wire42(18);
	sub_wire1(22, 19)    <= sub_wire42(19);
	sub_wire1(22, 20)    <= sub_wire42(20);
	sub_wire1(22, 21)    <= sub_wire42(21);
	sub_wire1(22, 22)    <= sub_wire42(22);
	sub_wire1(22, 23)    <= sub_wire42(23);
	sub_wire1(22, 24)    <= sub_wire42(24);
	sub_wire1(22, 25)    <= sub_wire42(25);
	sub_wire1(22, 26)    <= sub_wire42(26);
	sub_wire1(22, 27)    <= sub_wire42(27);
	sub_wire1(22, 28)    <= sub_wire42(28);
	sub_wire1(22, 29)    <= sub_wire42(29);
	sub_wire1(22, 30)    <= sub_wire42(30);
	sub_wire1(22, 31)    <= sub_wire42(31);
	sub_wire1(21, 0)    <= sub_wire43(0);
	sub_wire1(21, 1)    <= sub_wire43(1);
	sub_wire1(21, 2)    <= sub_wire43(2);
	sub_wire1(21, 3)    <= sub_wire43(3);
	sub_wire1(21, 4)    <= sub_wire43(4);
	sub_wire1(21, 5)    <= sub_wire43(5);
	sub_wire1(21, 6)    <= sub_wire43(6);
	sub_wire1(21, 7)    <= sub_wire43(7);
	sub_wire1(21, 8)    <= sub_wire43(8);
	sub_wire1(21, 9)    <= sub_wire43(9);
	sub_wire1(21, 10)    <= sub_wire43(10);
	sub_wire1(21, 11)    <= sub_wire43(11);
	sub_wire1(21, 12)    <= sub_wire43(12);
	sub_wire1(21, 13)    <= sub_wire43(13);
	sub_wire1(21, 14)    <= sub_wire43(14);
	sub_wire1(21, 15)    <= sub_wire43(15);
	sub_wire1(21, 16)    <= sub_wire43(16);
	sub_wire1(21, 17)    <= sub_wire43(17);
	sub_wire1(21, 18)    <= sub_wire43(18);
	sub_wire1(21, 19)    <= sub_wire43(19);
	sub_wire1(21, 20)    <= sub_wire43(20);
	sub_wire1(21, 21)    <= sub_wire43(21);
	sub_wire1(21, 22)    <= sub_wire43(22);
	sub_wire1(21, 23)    <= sub_wire43(23);
	sub_wire1(21, 24)    <= sub_wire43(24);
	sub_wire1(21, 25)    <= sub_wire43(25);
	sub_wire1(21, 26)    <= sub_wire43(26);
	sub_wire1(21, 27)    <= sub_wire43(27);
	sub_wire1(21, 28)    <= sub_wire43(28);
	sub_wire1(21, 29)    <= sub_wire43(29);
	sub_wire1(21, 30)    <= sub_wire43(30);
	sub_wire1(21, 31)    <= sub_wire43(31);
	sub_wire1(20, 0)    <= sub_wire44(0);
	sub_wire1(20, 1)    <= sub_wire44(1);
	sub_wire1(20, 2)    <= sub_wire44(2);
	sub_wire1(20, 3)    <= sub_wire44(3);
	sub_wire1(20, 4)    <= sub_wire44(4);
	sub_wire1(20, 5)    <= sub_wire44(5);
	sub_wire1(20, 6)    <= sub_wire44(6);
	sub_wire1(20, 7)    <= sub_wire44(7);
	sub_wire1(20, 8)    <= sub_wire44(8);
	sub_wire1(20, 9)    <= sub_wire44(9);
	sub_wire1(20, 10)    <= sub_wire44(10);
	sub_wire1(20, 11)    <= sub_wire44(11);
	sub_wire1(20, 12)    <= sub_wire44(12);
	sub_wire1(20, 13)    <= sub_wire44(13);
	sub_wire1(20, 14)    <= sub_wire44(14);
	sub_wire1(20, 15)    <= sub_wire44(15);
	sub_wire1(20, 16)    <= sub_wire44(16);
	sub_wire1(20, 17)    <= sub_wire44(17);
	sub_wire1(20, 18)    <= sub_wire44(18);
	sub_wire1(20, 19)    <= sub_wire44(19);
	sub_wire1(20, 20)    <= sub_wire44(20);
	sub_wire1(20, 21)    <= sub_wire44(21);
	sub_wire1(20, 22)    <= sub_wire44(22);
	sub_wire1(20, 23)    <= sub_wire44(23);
	sub_wire1(20, 24)    <= sub_wire44(24);
	sub_wire1(20, 25)    <= sub_wire44(25);
	sub_wire1(20, 26)    <= sub_wire44(26);
	sub_wire1(20, 27)    <= sub_wire44(27);
	sub_wire1(20, 28)    <= sub_wire44(28);
	sub_wire1(20, 29)    <= sub_wire44(29);
	sub_wire1(20, 30)    <= sub_wire44(30);
	sub_wire1(20, 31)    <= sub_wire44(31);
	sub_wire1(19, 0)    <= sub_wire45(0);
	sub_wire1(19, 1)    <= sub_wire45(1);
	sub_wire1(19, 2)    <= sub_wire45(2);
	sub_wire1(19, 3)    <= sub_wire45(3);
	sub_wire1(19, 4)    <= sub_wire45(4);
	sub_wire1(19, 5)    <= sub_wire45(5);
	sub_wire1(19, 6)    <= sub_wire45(6);
	sub_wire1(19, 7)    <= sub_wire45(7);
	sub_wire1(19, 8)    <= sub_wire45(8);
	sub_wire1(19, 9)    <= sub_wire45(9);
	sub_wire1(19, 10)    <= sub_wire45(10);
	sub_wire1(19, 11)    <= sub_wire45(11);
	sub_wire1(19, 12)    <= sub_wire45(12);
	sub_wire1(19, 13)    <= sub_wire45(13);
	sub_wire1(19, 14)    <= sub_wire45(14);
	sub_wire1(19, 15)    <= sub_wire45(15);
	sub_wire1(19, 16)    <= sub_wire45(16);
	sub_wire1(19, 17)    <= sub_wire45(17);
	sub_wire1(19, 18)    <= sub_wire45(18);
	sub_wire1(19, 19)    <= sub_wire45(19);
	sub_wire1(19, 20)    <= sub_wire45(20);
	sub_wire1(19, 21)    <= sub_wire45(21);
	sub_wire1(19, 22)    <= sub_wire45(22);
	sub_wire1(19, 23)    <= sub_wire45(23);
	sub_wire1(19, 24)    <= sub_wire45(24);
	sub_wire1(19, 25)    <= sub_wire45(25);
	sub_wire1(19, 26)    <= sub_wire45(26);
	sub_wire1(19, 27)    <= sub_wire45(27);
	sub_wire1(19, 28)    <= sub_wire45(28);
	sub_wire1(19, 29)    <= sub_wire45(29);
	sub_wire1(19, 30)    <= sub_wire45(30);
	sub_wire1(19, 31)    <= sub_wire45(31);
	sub_wire1(18, 0)    <= sub_wire46(0);
	sub_wire1(18, 1)    <= sub_wire46(1);
	sub_wire1(18, 2)    <= sub_wire46(2);
	sub_wire1(18, 3)    <= sub_wire46(3);
	sub_wire1(18, 4)    <= sub_wire46(4);
	sub_wire1(18, 5)    <= sub_wire46(5);
	sub_wire1(18, 6)    <= sub_wire46(6);
	sub_wire1(18, 7)    <= sub_wire46(7);
	sub_wire1(18, 8)    <= sub_wire46(8);
	sub_wire1(18, 9)    <= sub_wire46(9);
	sub_wire1(18, 10)    <= sub_wire46(10);
	sub_wire1(18, 11)    <= sub_wire46(11);
	sub_wire1(18, 12)    <= sub_wire46(12);
	sub_wire1(18, 13)    <= sub_wire46(13);
	sub_wire1(18, 14)    <= sub_wire46(14);
	sub_wire1(18, 15)    <= sub_wire46(15);
	sub_wire1(18, 16)    <= sub_wire46(16);
	sub_wire1(18, 17)    <= sub_wire46(17);
	sub_wire1(18, 18)    <= sub_wire46(18);
	sub_wire1(18, 19)    <= sub_wire46(19);
	sub_wire1(18, 20)    <= sub_wire46(20);
	sub_wire1(18, 21)    <= sub_wire46(21);
	sub_wire1(18, 22)    <= sub_wire46(22);
	sub_wire1(18, 23)    <= sub_wire46(23);
	sub_wire1(18, 24)    <= sub_wire46(24);
	sub_wire1(18, 25)    <= sub_wire46(25);
	sub_wire1(18, 26)    <= sub_wire46(26);
	sub_wire1(18, 27)    <= sub_wire46(27);
	sub_wire1(18, 28)    <= sub_wire46(28);
	sub_wire1(18, 29)    <= sub_wire46(29);
	sub_wire1(18, 30)    <= sub_wire46(30);
	sub_wire1(18, 31)    <= sub_wire46(31);
	sub_wire1(17, 0)    <= sub_wire47(0);
	sub_wire1(17, 1)    <= sub_wire47(1);
	sub_wire1(17, 2)    <= sub_wire47(2);
	sub_wire1(17, 3)    <= sub_wire47(3);
	sub_wire1(17, 4)    <= sub_wire47(4);
	sub_wire1(17, 5)    <= sub_wire47(5);
	sub_wire1(17, 6)    <= sub_wire47(6);
	sub_wire1(17, 7)    <= sub_wire47(7);
	sub_wire1(17, 8)    <= sub_wire47(8);
	sub_wire1(17, 9)    <= sub_wire47(9);
	sub_wire1(17, 10)    <= sub_wire47(10);
	sub_wire1(17, 11)    <= sub_wire47(11);
	sub_wire1(17, 12)    <= sub_wire47(12);
	sub_wire1(17, 13)    <= sub_wire47(13);
	sub_wire1(17, 14)    <= sub_wire47(14);
	sub_wire1(17, 15)    <= sub_wire47(15);
	sub_wire1(17, 16)    <= sub_wire47(16);
	sub_wire1(17, 17)    <= sub_wire47(17);
	sub_wire1(17, 18)    <= sub_wire47(18);
	sub_wire1(17, 19)    <= sub_wire47(19);
	sub_wire1(17, 20)    <= sub_wire47(20);
	sub_wire1(17, 21)    <= sub_wire47(21);
	sub_wire1(17, 22)    <= sub_wire47(22);
	sub_wire1(17, 23)    <= sub_wire47(23);
	sub_wire1(17, 24)    <= sub_wire47(24);
	sub_wire1(17, 25)    <= sub_wire47(25);
	sub_wire1(17, 26)    <= sub_wire47(26);
	sub_wire1(17, 27)    <= sub_wire47(27);
	sub_wire1(17, 28)    <= sub_wire47(28);
	sub_wire1(17, 29)    <= sub_wire47(29);
	sub_wire1(17, 30)    <= sub_wire47(30);
	sub_wire1(17, 31)    <= sub_wire47(31);
	sub_wire1(16, 0)    <= sub_wire48(0);
	sub_wire1(16, 1)    <= sub_wire48(1);
	sub_wire1(16, 2)    <= sub_wire48(2);
	sub_wire1(16, 3)    <= sub_wire48(3);
	sub_wire1(16, 4)    <= sub_wire48(4);
	sub_wire1(16, 5)    <= sub_wire48(5);
	sub_wire1(16, 6)    <= sub_wire48(6);
	sub_wire1(16, 7)    <= sub_wire48(7);
	sub_wire1(16, 8)    <= sub_wire48(8);
	sub_wire1(16, 9)    <= sub_wire48(9);
	sub_wire1(16, 10)    <= sub_wire48(10);
	sub_wire1(16, 11)    <= sub_wire48(11);
	sub_wire1(16, 12)    <= sub_wire48(12);
	sub_wire1(16, 13)    <= sub_wire48(13);
	sub_wire1(16, 14)    <= sub_wire48(14);
	sub_wire1(16, 15)    <= sub_wire48(15);
	sub_wire1(16, 16)    <= sub_wire48(16);
	sub_wire1(16, 17)    <= sub_wire48(17);
	sub_wire1(16, 18)    <= sub_wire48(18);
	sub_wire1(16, 19)    <= sub_wire48(19);
	sub_wire1(16, 20)    <= sub_wire48(20);
	sub_wire1(16, 21)    <= sub_wire48(21);
	sub_wire1(16, 22)    <= sub_wire48(22);
	sub_wire1(16, 23)    <= sub_wire48(23);
	sub_wire1(16, 24)    <= sub_wire48(24);
	sub_wire1(16, 25)    <= sub_wire48(25);
	sub_wire1(16, 26)    <= sub_wire48(26);
	sub_wire1(16, 27)    <= sub_wire48(27);
	sub_wire1(16, 28)    <= sub_wire48(28);
	sub_wire1(16, 29)    <= sub_wire48(29);
	sub_wire1(16, 30)    <= sub_wire48(30);
	sub_wire1(16, 31)    <= sub_wire48(31);
	sub_wire1(15, 0)    <= sub_wire49(0);
	sub_wire1(15, 1)    <= sub_wire49(1);
	sub_wire1(15, 2)    <= sub_wire49(2);
	sub_wire1(15, 3)    <= sub_wire49(3);
	sub_wire1(15, 4)    <= sub_wire49(4);
	sub_wire1(15, 5)    <= sub_wire49(5);
	sub_wire1(15, 6)    <= sub_wire49(6);
	sub_wire1(15, 7)    <= sub_wire49(7);
	sub_wire1(15, 8)    <= sub_wire49(8);
	sub_wire1(15, 9)    <= sub_wire49(9);
	sub_wire1(15, 10)    <= sub_wire49(10);
	sub_wire1(15, 11)    <= sub_wire49(11);
	sub_wire1(15, 12)    <= sub_wire49(12);
	sub_wire1(15, 13)    <= sub_wire49(13);
	sub_wire1(15, 14)    <= sub_wire49(14);
	sub_wire1(15, 15)    <= sub_wire49(15);
	sub_wire1(15, 16)    <= sub_wire49(16);
	sub_wire1(15, 17)    <= sub_wire49(17);
	sub_wire1(15, 18)    <= sub_wire49(18);
	sub_wire1(15, 19)    <= sub_wire49(19);
	sub_wire1(15, 20)    <= sub_wire49(20);
	sub_wire1(15, 21)    <= sub_wire49(21);
	sub_wire1(15, 22)    <= sub_wire49(22);
	sub_wire1(15, 23)    <= sub_wire49(23);
	sub_wire1(15, 24)    <= sub_wire49(24);
	sub_wire1(15, 25)    <= sub_wire49(25);
	sub_wire1(15, 26)    <= sub_wire49(26);
	sub_wire1(15, 27)    <= sub_wire49(27);
	sub_wire1(15, 28)    <= sub_wire49(28);
	sub_wire1(15, 29)    <= sub_wire49(29);
	sub_wire1(15, 30)    <= sub_wire49(30);
	sub_wire1(15, 31)    <= sub_wire49(31);
	sub_wire1(14, 0)    <= sub_wire50(0);
	sub_wire1(14, 1)    <= sub_wire50(1);
	sub_wire1(14, 2)    <= sub_wire50(2);
	sub_wire1(14, 3)    <= sub_wire50(3);
	sub_wire1(14, 4)    <= sub_wire50(4);
	sub_wire1(14, 5)    <= sub_wire50(5);
	sub_wire1(14, 6)    <= sub_wire50(6);
	sub_wire1(14, 7)    <= sub_wire50(7);
	sub_wire1(14, 8)    <= sub_wire50(8);
	sub_wire1(14, 9)    <= sub_wire50(9);
	sub_wire1(14, 10)    <= sub_wire50(10);
	sub_wire1(14, 11)    <= sub_wire50(11);
	sub_wire1(14, 12)    <= sub_wire50(12);
	sub_wire1(14, 13)    <= sub_wire50(13);
	sub_wire1(14, 14)    <= sub_wire50(14);
	sub_wire1(14, 15)    <= sub_wire50(15);
	sub_wire1(14, 16)    <= sub_wire50(16);
	sub_wire1(14, 17)    <= sub_wire50(17);
	sub_wire1(14, 18)    <= sub_wire50(18);
	sub_wire1(14, 19)    <= sub_wire50(19);
	sub_wire1(14, 20)    <= sub_wire50(20);
	sub_wire1(14, 21)    <= sub_wire50(21);
	sub_wire1(14, 22)    <= sub_wire50(22);
	sub_wire1(14, 23)    <= sub_wire50(23);
	sub_wire1(14, 24)    <= sub_wire50(24);
	sub_wire1(14, 25)    <= sub_wire50(25);
	sub_wire1(14, 26)    <= sub_wire50(26);
	sub_wire1(14, 27)    <= sub_wire50(27);
	sub_wire1(14, 28)    <= sub_wire50(28);
	sub_wire1(14, 29)    <= sub_wire50(29);
	sub_wire1(14, 30)    <= sub_wire50(30);
	sub_wire1(14, 31)    <= sub_wire50(31);
	sub_wire1(13, 0)    <= sub_wire51(0);
	sub_wire1(13, 1)    <= sub_wire51(1);
	sub_wire1(13, 2)    <= sub_wire51(2);
	sub_wire1(13, 3)    <= sub_wire51(3);
	sub_wire1(13, 4)    <= sub_wire51(4);
	sub_wire1(13, 5)    <= sub_wire51(5);
	sub_wire1(13, 6)    <= sub_wire51(6);
	sub_wire1(13, 7)    <= sub_wire51(7);
	sub_wire1(13, 8)    <= sub_wire51(8);
	sub_wire1(13, 9)    <= sub_wire51(9);
	sub_wire1(13, 10)    <= sub_wire51(10);
	sub_wire1(13, 11)    <= sub_wire51(11);
	sub_wire1(13, 12)    <= sub_wire51(12);
	sub_wire1(13, 13)    <= sub_wire51(13);
	sub_wire1(13, 14)    <= sub_wire51(14);
	sub_wire1(13, 15)    <= sub_wire51(15);
	sub_wire1(13, 16)    <= sub_wire51(16);
	sub_wire1(13, 17)    <= sub_wire51(17);
	sub_wire1(13, 18)    <= sub_wire51(18);
	sub_wire1(13, 19)    <= sub_wire51(19);
	sub_wire1(13, 20)    <= sub_wire51(20);
	sub_wire1(13, 21)    <= sub_wire51(21);
	sub_wire1(13, 22)    <= sub_wire51(22);
	sub_wire1(13, 23)    <= sub_wire51(23);
	sub_wire1(13, 24)    <= sub_wire51(24);
	sub_wire1(13, 25)    <= sub_wire51(25);
	sub_wire1(13, 26)    <= sub_wire51(26);
	sub_wire1(13, 27)    <= sub_wire51(27);
	sub_wire1(13, 28)    <= sub_wire51(28);
	sub_wire1(13, 29)    <= sub_wire51(29);
	sub_wire1(13, 30)    <= sub_wire51(30);
	sub_wire1(13, 31)    <= sub_wire51(31);
	sub_wire1(12, 0)    <= sub_wire52(0);
	sub_wire1(12, 1)    <= sub_wire52(1);
	sub_wire1(12, 2)    <= sub_wire52(2);
	sub_wire1(12, 3)    <= sub_wire52(3);
	sub_wire1(12, 4)    <= sub_wire52(4);
	sub_wire1(12, 5)    <= sub_wire52(5);
	sub_wire1(12, 6)    <= sub_wire52(6);
	sub_wire1(12, 7)    <= sub_wire52(7);
	sub_wire1(12, 8)    <= sub_wire52(8);
	sub_wire1(12, 9)    <= sub_wire52(9);
	sub_wire1(12, 10)    <= sub_wire52(10);
	sub_wire1(12, 11)    <= sub_wire52(11);
	sub_wire1(12, 12)    <= sub_wire52(12);
	sub_wire1(12, 13)    <= sub_wire52(13);
	sub_wire1(12, 14)    <= sub_wire52(14);
	sub_wire1(12, 15)    <= sub_wire52(15);
	sub_wire1(12, 16)    <= sub_wire52(16);
	sub_wire1(12, 17)    <= sub_wire52(17);
	sub_wire1(12, 18)    <= sub_wire52(18);
	sub_wire1(12, 19)    <= sub_wire52(19);
	sub_wire1(12, 20)    <= sub_wire52(20);
	sub_wire1(12, 21)    <= sub_wire52(21);
	sub_wire1(12, 22)    <= sub_wire52(22);
	sub_wire1(12, 23)    <= sub_wire52(23);
	sub_wire1(12, 24)    <= sub_wire52(24);
	sub_wire1(12, 25)    <= sub_wire52(25);
	sub_wire1(12, 26)    <= sub_wire52(26);
	sub_wire1(12, 27)    <= sub_wire52(27);
	sub_wire1(12, 28)    <= sub_wire52(28);
	sub_wire1(12, 29)    <= sub_wire52(29);
	sub_wire1(12, 30)    <= sub_wire52(30);
	sub_wire1(12, 31)    <= sub_wire52(31);
	sub_wire1(11, 0)    <= sub_wire53(0);
	sub_wire1(11, 1)    <= sub_wire53(1);
	sub_wire1(11, 2)    <= sub_wire53(2);
	sub_wire1(11, 3)    <= sub_wire53(3);
	sub_wire1(11, 4)    <= sub_wire53(4);
	sub_wire1(11, 5)    <= sub_wire53(5);
	sub_wire1(11, 6)    <= sub_wire53(6);
	sub_wire1(11, 7)    <= sub_wire53(7);
	sub_wire1(11, 8)    <= sub_wire53(8);
	sub_wire1(11, 9)    <= sub_wire53(9);
	sub_wire1(11, 10)    <= sub_wire53(10);
	sub_wire1(11, 11)    <= sub_wire53(11);
	sub_wire1(11, 12)    <= sub_wire53(12);
	sub_wire1(11, 13)    <= sub_wire53(13);
	sub_wire1(11, 14)    <= sub_wire53(14);
	sub_wire1(11, 15)    <= sub_wire53(15);
	sub_wire1(11, 16)    <= sub_wire53(16);
	sub_wire1(11, 17)    <= sub_wire53(17);
	sub_wire1(11, 18)    <= sub_wire53(18);
	sub_wire1(11, 19)    <= sub_wire53(19);
	sub_wire1(11, 20)    <= sub_wire53(20);
	sub_wire1(11, 21)    <= sub_wire53(21);
	sub_wire1(11, 22)    <= sub_wire53(22);
	sub_wire1(11, 23)    <= sub_wire53(23);
	sub_wire1(11, 24)    <= sub_wire53(24);
	sub_wire1(11, 25)    <= sub_wire53(25);
	sub_wire1(11, 26)    <= sub_wire53(26);
	sub_wire1(11, 27)    <= sub_wire53(27);
	sub_wire1(11, 28)    <= sub_wire53(28);
	sub_wire1(11, 29)    <= sub_wire53(29);
	sub_wire1(11, 30)    <= sub_wire53(30);
	sub_wire1(11, 31)    <= sub_wire53(31);
	sub_wire1(10, 0)    <= sub_wire54(0);
	sub_wire1(10, 1)    <= sub_wire54(1);
	sub_wire1(10, 2)    <= sub_wire54(2);
	sub_wire1(10, 3)    <= sub_wire54(3);
	sub_wire1(10, 4)    <= sub_wire54(4);
	sub_wire1(10, 5)    <= sub_wire54(5);
	sub_wire1(10, 6)    <= sub_wire54(6);
	sub_wire1(10, 7)    <= sub_wire54(7);
	sub_wire1(10, 8)    <= sub_wire54(8);
	sub_wire1(10, 9)    <= sub_wire54(9);
	sub_wire1(10, 10)    <= sub_wire54(10);
	sub_wire1(10, 11)    <= sub_wire54(11);
	sub_wire1(10, 12)    <= sub_wire54(12);
	sub_wire1(10, 13)    <= sub_wire54(13);
	sub_wire1(10, 14)    <= sub_wire54(14);
	sub_wire1(10, 15)    <= sub_wire54(15);
	sub_wire1(10, 16)    <= sub_wire54(16);
	sub_wire1(10, 17)    <= sub_wire54(17);
	sub_wire1(10, 18)    <= sub_wire54(18);
	sub_wire1(10, 19)    <= sub_wire54(19);
	sub_wire1(10, 20)    <= sub_wire54(20);
	sub_wire1(10, 21)    <= sub_wire54(21);
	sub_wire1(10, 22)    <= sub_wire54(22);
	sub_wire1(10, 23)    <= sub_wire54(23);
	sub_wire1(10, 24)    <= sub_wire54(24);
	sub_wire1(10, 25)    <= sub_wire54(25);
	sub_wire1(10, 26)    <= sub_wire54(26);
	sub_wire1(10, 27)    <= sub_wire54(27);
	sub_wire1(10, 28)    <= sub_wire54(28);
	sub_wire1(10, 29)    <= sub_wire54(29);
	sub_wire1(10, 30)    <= sub_wire54(30);
	sub_wire1(10, 31)    <= sub_wire54(31);
	sub_wire1(9, 0)    <= sub_wire55(0);
	sub_wire1(9, 1)    <= sub_wire55(1);
	sub_wire1(9, 2)    <= sub_wire55(2);
	sub_wire1(9, 3)    <= sub_wire55(3);
	sub_wire1(9, 4)    <= sub_wire55(4);
	sub_wire1(9, 5)    <= sub_wire55(5);
	sub_wire1(9, 6)    <= sub_wire55(6);
	sub_wire1(9, 7)    <= sub_wire55(7);
	sub_wire1(9, 8)    <= sub_wire55(8);
	sub_wire1(9, 9)    <= sub_wire55(9);
	sub_wire1(9, 10)    <= sub_wire55(10);
	sub_wire1(9, 11)    <= sub_wire55(11);
	sub_wire1(9, 12)    <= sub_wire55(12);
	sub_wire1(9, 13)    <= sub_wire55(13);
	sub_wire1(9, 14)    <= sub_wire55(14);
	sub_wire1(9, 15)    <= sub_wire55(15);
	sub_wire1(9, 16)    <= sub_wire55(16);
	sub_wire1(9, 17)    <= sub_wire55(17);
	sub_wire1(9, 18)    <= sub_wire55(18);
	sub_wire1(9, 19)    <= sub_wire55(19);
	sub_wire1(9, 20)    <= sub_wire55(20);
	sub_wire1(9, 21)    <= sub_wire55(21);
	sub_wire1(9, 22)    <= sub_wire55(22);
	sub_wire1(9, 23)    <= sub_wire55(23);
	sub_wire1(9, 24)    <= sub_wire55(24);
	sub_wire1(9, 25)    <= sub_wire55(25);
	sub_wire1(9, 26)    <= sub_wire55(26);
	sub_wire1(9, 27)    <= sub_wire55(27);
	sub_wire1(9, 28)    <= sub_wire55(28);
	sub_wire1(9, 29)    <= sub_wire55(29);
	sub_wire1(9, 30)    <= sub_wire55(30);
	sub_wire1(9, 31)    <= sub_wire55(31);
	sub_wire1(8, 0)    <= sub_wire56(0);
	sub_wire1(8, 1)    <= sub_wire56(1);
	sub_wire1(8, 2)    <= sub_wire56(2);
	sub_wire1(8, 3)    <= sub_wire56(3);
	sub_wire1(8, 4)    <= sub_wire56(4);
	sub_wire1(8, 5)    <= sub_wire56(5);
	sub_wire1(8, 6)    <= sub_wire56(6);
	sub_wire1(8, 7)    <= sub_wire56(7);
	sub_wire1(8, 8)    <= sub_wire56(8);
	sub_wire1(8, 9)    <= sub_wire56(9);
	sub_wire1(8, 10)    <= sub_wire56(10);
	sub_wire1(8, 11)    <= sub_wire56(11);
	sub_wire1(8, 12)    <= sub_wire56(12);
	sub_wire1(8, 13)    <= sub_wire56(13);
	sub_wire1(8, 14)    <= sub_wire56(14);
	sub_wire1(8, 15)    <= sub_wire56(15);
	sub_wire1(8, 16)    <= sub_wire56(16);
	sub_wire1(8, 17)    <= sub_wire56(17);
	sub_wire1(8, 18)    <= sub_wire56(18);
	sub_wire1(8, 19)    <= sub_wire56(19);
	sub_wire1(8, 20)    <= sub_wire56(20);
	sub_wire1(8, 21)    <= sub_wire56(21);
	sub_wire1(8, 22)    <= sub_wire56(22);
	sub_wire1(8, 23)    <= sub_wire56(23);
	sub_wire1(8, 24)    <= sub_wire56(24);
	sub_wire1(8, 25)    <= sub_wire56(25);
	sub_wire1(8, 26)    <= sub_wire56(26);
	sub_wire1(8, 27)    <= sub_wire56(27);
	sub_wire1(8, 28)    <= sub_wire56(28);
	sub_wire1(8, 29)    <= sub_wire56(29);
	sub_wire1(8, 30)    <= sub_wire56(30);
	sub_wire1(8, 31)    <= sub_wire56(31);
	sub_wire1(7, 0)    <= sub_wire57(0);
	sub_wire1(7, 1)    <= sub_wire57(1);
	sub_wire1(7, 2)    <= sub_wire57(2);
	sub_wire1(7, 3)    <= sub_wire57(3);
	sub_wire1(7, 4)    <= sub_wire57(4);
	sub_wire1(7, 5)    <= sub_wire57(5);
	sub_wire1(7, 6)    <= sub_wire57(6);
	sub_wire1(7, 7)    <= sub_wire57(7);
	sub_wire1(7, 8)    <= sub_wire57(8);
	sub_wire1(7, 9)    <= sub_wire57(9);
	sub_wire1(7, 10)    <= sub_wire57(10);
	sub_wire1(7, 11)    <= sub_wire57(11);
	sub_wire1(7, 12)    <= sub_wire57(12);
	sub_wire1(7, 13)    <= sub_wire57(13);
	sub_wire1(7, 14)    <= sub_wire57(14);
	sub_wire1(7, 15)    <= sub_wire57(15);
	sub_wire1(7, 16)    <= sub_wire57(16);
	sub_wire1(7, 17)    <= sub_wire57(17);
	sub_wire1(7, 18)    <= sub_wire57(18);
	sub_wire1(7, 19)    <= sub_wire57(19);
	sub_wire1(7, 20)    <= sub_wire57(20);
	sub_wire1(7, 21)    <= sub_wire57(21);
	sub_wire1(7, 22)    <= sub_wire57(22);
	sub_wire1(7, 23)    <= sub_wire57(23);
	sub_wire1(7, 24)    <= sub_wire57(24);
	sub_wire1(7, 25)    <= sub_wire57(25);
	sub_wire1(7, 26)    <= sub_wire57(26);
	sub_wire1(7, 27)    <= sub_wire57(27);
	sub_wire1(7, 28)    <= sub_wire57(28);
	sub_wire1(7, 29)    <= sub_wire57(29);
	sub_wire1(7, 30)    <= sub_wire57(30);
	sub_wire1(7, 31)    <= sub_wire57(31);
	sub_wire1(6, 0)    <= sub_wire58(0);
	sub_wire1(6, 1)    <= sub_wire58(1);
	sub_wire1(6, 2)    <= sub_wire58(2);
	sub_wire1(6, 3)    <= sub_wire58(3);
	sub_wire1(6, 4)    <= sub_wire58(4);
	sub_wire1(6, 5)    <= sub_wire58(5);
	sub_wire1(6, 6)    <= sub_wire58(6);
	sub_wire1(6, 7)    <= sub_wire58(7);
	sub_wire1(6, 8)    <= sub_wire58(8);
	sub_wire1(6, 9)    <= sub_wire58(9);
	sub_wire1(6, 10)    <= sub_wire58(10);
	sub_wire1(6, 11)    <= sub_wire58(11);
	sub_wire1(6, 12)    <= sub_wire58(12);
	sub_wire1(6, 13)    <= sub_wire58(13);
	sub_wire1(6, 14)    <= sub_wire58(14);
	sub_wire1(6, 15)    <= sub_wire58(15);
	sub_wire1(6, 16)    <= sub_wire58(16);
	sub_wire1(6, 17)    <= sub_wire58(17);
	sub_wire1(6, 18)    <= sub_wire58(18);
	sub_wire1(6, 19)    <= sub_wire58(19);
	sub_wire1(6, 20)    <= sub_wire58(20);
	sub_wire1(6, 21)    <= sub_wire58(21);
	sub_wire1(6, 22)    <= sub_wire58(22);
	sub_wire1(6, 23)    <= sub_wire58(23);
	sub_wire1(6, 24)    <= sub_wire58(24);
	sub_wire1(6, 25)    <= sub_wire58(25);
	sub_wire1(6, 26)    <= sub_wire58(26);
	sub_wire1(6, 27)    <= sub_wire58(27);
	sub_wire1(6, 28)    <= sub_wire58(28);
	sub_wire1(6, 29)    <= sub_wire58(29);
	sub_wire1(6, 30)    <= sub_wire58(30);
	sub_wire1(6, 31)    <= sub_wire58(31);
	sub_wire1(5, 0)    <= sub_wire59(0);
	sub_wire1(5, 1)    <= sub_wire59(1);
	sub_wire1(5, 2)    <= sub_wire59(2);
	sub_wire1(5, 3)    <= sub_wire59(3);
	sub_wire1(5, 4)    <= sub_wire59(4);
	sub_wire1(5, 5)    <= sub_wire59(5);
	sub_wire1(5, 6)    <= sub_wire59(6);
	sub_wire1(5, 7)    <= sub_wire59(7);
	sub_wire1(5, 8)    <= sub_wire59(8);
	sub_wire1(5, 9)    <= sub_wire59(9);
	sub_wire1(5, 10)    <= sub_wire59(10);
	sub_wire1(5, 11)    <= sub_wire59(11);
	sub_wire1(5, 12)    <= sub_wire59(12);
	sub_wire1(5, 13)    <= sub_wire59(13);
	sub_wire1(5, 14)    <= sub_wire59(14);
	sub_wire1(5, 15)    <= sub_wire59(15);
	sub_wire1(5, 16)    <= sub_wire59(16);
	sub_wire1(5, 17)    <= sub_wire59(17);
	sub_wire1(5, 18)    <= sub_wire59(18);
	sub_wire1(5, 19)    <= sub_wire59(19);
	sub_wire1(5, 20)    <= sub_wire59(20);
	sub_wire1(5, 21)    <= sub_wire59(21);
	sub_wire1(5, 22)    <= sub_wire59(22);
	sub_wire1(5, 23)    <= sub_wire59(23);
	sub_wire1(5, 24)    <= sub_wire59(24);
	sub_wire1(5, 25)    <= sub_wire59(25);
	sub_wire1(5, 26)    <= sub_wire59(26);
	sub_wire1(5, 27)    <= sub_wire59(27);
	sub_wire1(5, 28)    <= sub_wire59(28);
	sub_wire1(5, 29)    <= sub_wire59(29);
	sub_wire1(5, 30)    <= sub_wire59(30);
	sub_wire1(5, 31)    <= sub_wire59(31);
	sub_wire1(4, 0)    <= sub_wire60(0);
	sub_wire1(4, 1)    <= sub_wire60(1);
	sub_wire1(4, 2)    <= sub_wire60(2);
	sub_wire1(4, 3)    <= sub_wire60(3);
	sub_wire1(4, 4)    <= sub_wire60(4);
	sub_wire1(4, 5)    <= sub_wire60(5);
	sub_wire1(4, 6)    <= sub_wire60(6);
	sub_wire1(4, 7)    <= sub_wire60(7);
	sub_wire1(4, 8)    <= sub_wire60(8);
	sub_wire1(4, 9)    <= sub_wire60(9);
	sub_wire1(4, 10)    <= sub_wire60(10);
	sub_wire1(4, 11)    <= sub_wire60(11);
	sub_wire1(4, 12)    <= sub_wire60(12);
	sub_wire1(4, 13)    <= sub_wire60(13);
	sub_wire1(4, 14)    <= sub_wire60(14);
	sub_wire1(4, 15)    <= sub_wire60(15);
	sub_wire1(4, 16)    <= sub_wire60(16);
	sub_wire1(4, 17)    <= sub_wire60(17);
	sub_wire1(4, 18)    <= sub_wire60(18);
	sub_wire1(4, 19)    <= sub_wire60(19);
	sub_wire1(4, 20)    <= sub_wire60(20);
	sub_wire1(4, 21)    <= sub_wire60(21);
	sub_wire1(4, 22)    <= sub_wire60(22);
	sub_wire1(4, 23)    <= sub_wire60(23);
	sub_wire1(4, 24)    <= sub_wire60(24);
	sub_wire1(4, 25)    <= sub_wire60(25);
	sub_wire1(4, 26)    <= sub_wire60(26);
	sub_wire1(4, 27)    <= sub_wire60(27);
	sub_wire1(4, 28)    <= sub_wire60(28);
	sub_wire1(4, 29)    <= sub_wire60(29);
	sub_wire1(4, 30)    <= sub_wire60(30);
	sub_wire1(4, 31)    <= sub_wire60(31);
	sub_wire1(3, 0)    <= sub_wire61(0);
	sub_wire1(3, 1)    <= sub_wire61(1);
	sub_wire1(3, 2)    <= sub_wire61(2);
	sub_wire1(3, 3)    <= sub_wire61(3);
	sub_wire1(3, 4)    <= sub_wire61(4);
	sub_wire1(3, 5)    <= sub_wire61(5);
	sub_wire1(3, 6)    <= sub_wire61(6);
	sub_wire1(3, 7)    <= sub_wire61(7);
	sub_wire1(3, 8)    <= sub_wire61(8);
	sub_wire1(3, 9)    <= sub_wire61(9);
	sub_wire1(3, 10)    <= sub_wire61(10);
	sub_wire1(3, 11)    <= sub_wire61(11);
	sub_wire1(3, 12)    <= sub_wire61(12);
	sub_wire1(3, 13)    <= sub_wire61(13);
	sub_wire1(3, 14)    <= sub_wire61(14);
	sub_wire1(3, 15)    <= sub_wire61(15);
	sub_wire1(3, 16)    <= sub_wire61(16);
	sub_wire1(3, 17)    <= sub_wire61(17);
	sub_wire1(3, 18)    <= sub_wire61(18);
	sub_wire1(3, 19)    <= sub_wire61(19);
	sub_wire1(3, 20)    <= sub_wire61(20);
	sub_wire1(3, 21)    <= sub_wire61(21);
	sub_wire1(3, 22)    <= sub_wire61(22);
	sub_wire1(3, 23)    <= sub_wire61(23);
	sub_wire1(3, 24)    <= sub_wire61(24);
	sub_wire1(3, 25)    <= sub_wire61(25);
	sub_wire1(3, 26)    <= sub_wire61(26);
	sub_wire1(3, 27)    <= sub_wire61(27);
	sub_wire1(3, 28)    <= sub_wire61(28);
	sub_wire1(3, 29)    <= sub_wire61(29);
	sub_wire1(3, 30)    <= sub_wire61(30);
	sub_wire1(3, 31)    <= sub_wire61(31);
	sub_wire1(2, 0)    <= sub_wire62(0);
	sub_wire1(2, 1)    <= sub_wire62(1);
	sub_wire1(2, 2)    <= sub_wire62(2);
	sub_wire1(2, 3)    <= sub_wire62(3);
	sub_wire1(2, 4)    <= sub_wire62(4);
	sub_wire1(2, 5)    <= sub_wire62(5);
	sub_wire1(2, 6)    <= sub_wire62(6);
	sub_wire1(2, 7)    <= sub_wire62(7);
	sub_wire1(2, 8)    <= sub_wire62(8);
	sub_wire1(2, 9)    <= sub_wire62(9);
	sub_wire1(2, 10)    <= sub_wire62(10);
	sub_wire1(2, 11)    <= sub_wire62(11);
	sub_wire1(2, 12)    <= sub_wire62(12);
	sub_wire1(2, 13)    <= sub_wire62(13);
	sub_wire1(2, 14)    <= sub_wire62(14);
	sub_wire1(2, 15)    <= sub_wire62(15);
	sub_wire1(2, 16)    <= sub_wire62(16);
	sub_wire1(2, 17)    <= sub_wire62(17);
	sub_wire1(2, 18)    <= sub_wire62(18);
	sub_wire1(2, 19)    <= sub_wire62(19);
	sub_wire1(2, 20)    <= sub_wire62(20);
	sub_wire1(2, 21)    <= sub_wire62(21);
	sub_wire1(2, 22)    <= sub_wire62(22);
	sub_wire1(2, 23)    <= sub_wire62(23);
	sub_wire1(2, 24)    <= sub_wire62(24);
	sub_wire1(2, 25)    <= sub_wire62(25);
	sub_wire1(2, 26)    <= sub_wire62(26);
	sub_wire1(2, 27)    <= sub_wire62(27);
	sub_wire1(2, 28)    <= sub_wire62(28);
	sub_wire1(2, 29)    <= sub_wire62(29);
	sub_wire1(2, 30)    <= sub_wire62(30);
	sub_wire1(2, 31)    <= sub_wire62(31);
	sub_wire1(1, 0)    <= sub_wire63(0);
	sub_wire1(1, 1)    <= sub_wire63(1);
	sub_wire1(1, 2)    <= sub_wire63(2);
	sub_wire1(1, 3)    <= sub_wire63(3);
	sub_wire1(1, 4)    <= sub_wire63(4);
	sub_wire1(1, 5)    <= sub_wire63(5);
	sub_wire1(1, 6)    <= sub_wire63(6);
	sub_wire1(1, 7)    <= sub_wire63(7);
	sub_wire1(1, 8)    <= sub_wire63(8);
	sub_wire1(1, 9)    <= sub_wire63(9);
	sub_wire1(1, 10)    <= sub_wire63(10);
	sub_wire1(1, 11)    <= sub_wire63(11);
	sub_wire1(1, 12)    <= sub_wire63(12);
	sub_wire1(1, 13)    <= sub_wire63(13);
	sub_wire1(1, 14)    <= sub_wire63(14);
	sub_wire1(1, 15)    <= sub_wire63(15);
	sub_wire1(1, 16)    <= sub_wire63(16);
	sub_wire1(1, 17)    <= sub_wire63(17);
	sub_wire1(1, 18)    <= sub_wire63(18);
	sub_wire1(1, 19)    <= sub_wire63(19);
	sub_wire1(1, 20)    <= sub_wire63(20);
	sub_wire1(1, 21)    <= sub_wire63(21);
	sub_wire1(1, 22)    <= sub_wire63(22);
	sub_wire1(1, 23)    <= sub_wire63(23);
	sub_wire1(1, 24)    <= sub_wire63(24);
	sub_wire1(1, 25)    <= sub_wire63(25);
	sub_wire1(1, 26)    <= sub_wire63(26);
	sub_wire1(1, 27)    <= sub_wire63(27);
	sub_wire1(1, 28)    <= sub_wire63(28);
	sub_wire1(1, 29)    <= sub_wire63(29);
	sub_wire1(1, 30)    <= sub_wire63(30);
	sub_wire1(1, 31)    <= sub_wire63(31);
	sub_wire1(0, 0)    <= sub_wire64(0);
	sub_wire1(0, 1)    <= sub_wire64(1);
	sub_wire1(0, 2)    <= sub_wire64(2);
	sub_wire1(0, 3)    <= sub_wire64(3);
	sub_wire1(0, 4)    <= sub_wire64(4);
	sub_wire1(0, 5)    <= sub_wire64(5);
	sub_wire1(0, 6)    <= sub_wire64(6);
	sub_wire1(0, 7)    <= sub_wire64(7);
	sub_wire1(0, 8)    <= sub_wire64(8);
	sub_wire1(0, 9)    <= sub_wire64(9);
	sub_wire1(0, 10)    <= sub_wire64(10);
	sub_wire1(0, 11)    <= sub_wire64(11);
	sub_wire1(0, 12)    <= sub_wire64(12);
	sub_wire1(0, 13)    <= sub_wire64(13);
	sub_wire1(0, 14)    <= sub_wire64(14);
	sub_wire1(0, 15)    <= sub_wire64(15);
	sub_wire1(0, 16)    <= sub_wire64(16);
	sub_wire1(0, 17)    <= sub_wire64(17);
	sub_wire1(0, 18)    <= sub_wire64(18);
	sub_wire1(0, 19)    <= sub_wire64(19);
	sub_wire1(0, 20)    <= sub_wire64(20);
	sub_wire1(0, 21)    <= sub_wire64(21);
	sub_wire1(0, 22)    <= sub_wire64(22);
	sub_wire1(0, 23)    <= sub_wire64(23);
	sub_wire1(0, 24)    <= sub_wire64(24);
	sub_wire1(0, 25)    <= sub_wire64(25);
	sub_wire1(0, 26)    <= sub_wire64(26);
	sub_wire1(0, 27)    <= sub_wire64(27);
	sub_wire1(0, 28)    <= sub_wire64(28);
	sub_wire1(0, 29)    <= sub_wire64(29);
	sub_wire1(0, 30)    <= sub_wire64(30);
	sub_wire1(0, 31)    <= sub_wire64(31);
	result    <= sub_wire65(31 DOWNTO 0);

	LPM_MUX_component : LPM_MUX
	GENERIC MAP (
		lpm_size => 64,
		lpm_type => "LPM_MUX",
		lpm_width => 32,
		lpm_widths => 6
	)
	PORT MAP (
		data => sub_wire1,
		sel => sel,
		result => sub_wire65
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "64"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "32"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "6"
-- Retrieval info: USED_PORT: data0x 0 0 32 0 INPUT NODEFVAL "data0x[31..0]"
-- Retrieval info: USED_PORT: data10x 0 0 32 0 INPUT NODEFVAL "data10x[31..0]"
-- Retrieval info: USED_PORT: data11x 0 0 32 0 INPUT NODEFVAL "data11x[31..0]"
-- Retrieval info: USED_PORT: data12x 0 0 32 0 INPUT NODEFVAL "data12x[31..0]"
-- Retrieval info: USED_PORT: data13x 0 0 32 0 INPUT NODEFVAL "data13x[31..0]"
-- Retrieval info: USED_PORT: data14x 0 0 32 0 INPUT NODEFVAL "data14x[31..0]"
-- Retrieval info: USED_PORT: data15x 0 0 32 0 INPUT NODEFVAL "data15x[31..0]"
-- Retrieval info: USED_PORT: data16x 0 0 32 0 INPUT NODEFVAL "data16x[31..0]"
-- Retrieval info: USED_PORT: data17x 0 0 32 0 INPUT NODEFVAL "data17x[31..0]"
-- Retrieval info: USED_PORT: data18x 0 0 32 0 INPUT NODEFVAL "data18x[31..0]"
-- Retrieval info: USED_PORT: data19x 0 0 32 0 INPUT NODEFVAL "data19x[31..0]"
-- Retrieval info: USED_PORT: data1x 0 0 32 0 INPUT NODEFVAL "data1x[31..0]"
-- Retrieval info: USED_PORT: data20x 0 0 32 0 INPUT NODEFVAL "data20x[31..0]"
-- Retrieval info: USED_PORT: data21x 0 0 32 0 INPUT NODEFVAL "data21x[31..0]"
-- Retrieval info: USED_PORT: data22x 0 0 32 0 INPUT NODEFVAL "data22x[31..0]"
-- Retrieval info: USED_PORT: data23x 0 0 32 0 INPUT NODEFVAL "data23x[31..0]"
-- Retrieval info: USED_PORT: data24x 0 0 32 0 INPUT NODEFVAL "data24x[31..0]"
-- Retrieval info: USED_PORT: data25x 0 0 32 0 INPUT NODEFVAL "data25x[31..0]"
-- Retrieval info: USED_PORT: data26x 0 0 32 0 INPUT NODEFVAL "data26x[31..0]"
-- Retrieval info: USED_PORT: data27x 0 0 32 0 INPUT NODEFVAL "data27x[31..0]"
-- Retrieval info: USED_PORT: data28x 0 0 32 0 INPUT NODEFVAL "data28x[31..0]"
-- Retrieval info: USED_PORT: data29x 0 0 32 0 INPUT NODEFVAL "data29x[31..0]"
-- Retrieval info: USED_PORT: data2x 0 0 32 0 INPUT NODEFVAL "data2x[31..0]"
-- Retrieval info: USED_PORT: data30x 0 0 32 0 INPUT NODEFVAL "data30x[31..0]"
-- Retrieval info: USED_PORT: data31x 0 0 32 0 INPUT NODEFVAL "data31x[31..0]"
-- Retrieval info: USED_PORT: data32x 0 0 32 0 INPUT NODEFVAL "data32x[31..0]"
-- Retrieval info: USED_PORT: data33x 0 0 32 0 INPUT NODEFVAL "data33x[31..0]"
-- Retrieval info: USED_PORT: data34x 0 0 32 0 INPUT NODEFVAL "data34x[31..0]"
-- Retrieval info: USED_PORT: data35x 0 0 32 0 INPUT NODEFVAL "data35x[31..0]"
-- Retrieval info: USED_PORT: data36x 0 0 32 0 INPUT NODEFVAL "data36x[31..0]"
-- Retrieval info: USED_PORT: data37x 0 0 32 0 INPUT NODEFVAL "data37x[31..0]"
-- Retrieval info: USED_PORT: data38x 0 0 32 0 INPUT NODEFVAL "data38x[31..0]"
-- Retrieval info: USED_PORT: data39x 0 0 32 0 INPUT NODEFVAL "data39x[31..0]"
-- Retrieval info: USED_PORT: data3x 0 0 32 0 INPUT NODEFVAL "data3x[31..0]"
-- Retrieval info: USED_PORT: data40x 0 0 32 0 INPUT NODEFVAL "data40x[31..0]"
-- Retrieval info: USED_PORT: data41x 0 0 32 0 INPUT NODEFVAL "data41x[31..0]"
-- Retrieval info: USED_PORT: data42x 0 0 32 0 INPUT NODEFVAL "data42x[31..0]"
-- Retrieval info: USED_PORT: data43x 0 0 32 0 INPUT NODEFVAL "data43x[31..0]"
-- Retrieval info: USED_PORT: data44x 0 0 32 0 INPUT NODEFVAL "data44x[31..0]"
-- Retrieval info: USED_PORT: data45x 0 0 32 0 INPUT NODEFVAL "data45x[31..0]"
-- Retrieval info: USED_PORT: data46x 0 0 32 0 INPUT NODEFVAL "data46x[31..0]"
-- Retrieval info: USED_PORT: data47x 0 0 32 0 INPUT NODEFVAL "data47x[31..0]"
-- Retrieval info: USED_PORT: data48x 0 0 32 0 INPUT NODEFVAL "data48x[31..0]"
-- Retrieval info: USED_PORT: data49x 0 0 32 0 INPUT NODEFVAL "data49x[31..0]"
-- Retrieval info: USED_PORT: data4x 0 0 32 0 INPUT NODEFVAL "data4x[31..0]"
-- Retrieval info: USED_PORT: data50x 0 0 32 0 INPUT NODEFVAL "data50x[31..0]"
-- Retrieval info: USED_PORT: data51x 0 0 32 0 INPUT NODEFVAL "data51x[31..0]"
-- Retrieval info: USED_PORT: data52x 0 0 32 0 INPUT NODEFVAL "data52x[31..0]"
-- Retrieval info: USED_PORT: data53x 0 0 32 0 INPUT NODEFVAL "data53x[31..0]"
-- Retrieval info: USED_PORT: data54x 0 0 32 0 INPUT NODEFVAL "data54x[31..0]"
-- Retrieval info: USED_PORT: data55x 0 0 32 0 INPUT NODEFVAL "data55x[31..0]"
-- Retrieval info: USED_PORT: data56x 0 0 32 0 INPUT NODEFVAL "data56x[31..0]"
-- Retrieval info: USED_PORT: data57x 0 0 32 0 INPUT NODEFVAL "data57x[31..0]"
-- Retrieval info: USED_PORT: data58x 0 0 32 0 INPUT NODEFVAL "data58x[31..0]"
-- Retrieval info: USED_PORT: data59x 0 0 32 0 INPUT NODEFVAL "data59x[31..0]"
-- Retrieval info: USED_PORT: data5x 0 0 32 0 INPUT NODEFVAL "data5x[31..0]"
-- Retrieval info: USED_PORT: data60x 0 0 32 0 INPUT NODEFVAL "data60x[31..0]"
-- Retrieval info: USED_PORT: data61x 0 0 32 0 INPUT NODEFVAL "data61x[31..0]"
-- Retrieval info: USED_PORT: data62x 0 0 32 0 INPUT NODEFVAL "data62x[31..0]"
-- Retrieval info: USED_PORT: data63x 0 0 32 0 INPUT NODEFVAL "data63x[31..0]"
-- Retrieval info: USED_PORT: data6x 0 0 32 0 INPUT NODEFVAL "data6x[31..0]"
-- Retrieval info: USED_PORT: data7x 0 0 32 0 INPUT NODEFVAL "data7x[31..0]"
-- Retrieval info: USED_PORT: data8x 0 0 32 0 INPUT NODEFVAL "data8x[31..0]"
-- Retrieval info: USED_PORT: data9x 0 0 32 0 INPUT NODEFVAL "data9x[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: USED_PORT: sel 0 0 6 0 INPUT NODEFVAL "sel[5..0]"
-- Retrieval info: CONNECT: @data 1 0 32 0 data0x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 10 32 0 data10x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 11 32 0 data11x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 12 32 0 data12x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 13 32 0 data13x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 14 32 0 data14x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 15 32 0 data15x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 16 32 0 data16x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 17 32 0 data17x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 18 32 0 data18x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 19 32 0 data19x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 1 32 0 data1x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 20 32 0 data20x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 21 32 0 data21x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 22 32 0 data22x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 23 32 0 data23x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 24 32 0 data24x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 25 32 0 data25x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 26 32 0 data26x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 27 32 0 data27x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 28 32 0 data28x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 29 32 0 data29x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 2 32 0 data2x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 30 32 0 data30x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 31 32 0 data31x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 32 32 0 data32x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 33 32 0 data33x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 34 32 0 data34x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 35 32 0 data35x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 36 32 0 data36x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 37 32 0 data37x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 38 32 0 data38x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 39 32 0 data39x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 3 32 0 data3x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 40 32 0 data40x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 41 32 0 data41x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 42 32 0 data42x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 43 32 0 data43x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 44 32 0 data44x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 45 32 0 data45x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 46 32 0 data46x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 47 32 0 data47x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 48 32 0 data48x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 49 32 0 data49x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 4 32 0 data4x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 50 32 0 data50x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 51 32 0 data51x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 52 32 0 data52x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 53 32 0 data53x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 54 32 0 data54x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 55 32 0 data55x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 56 32 0 data56x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 57 32 0 data57x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 58 32 0 data58x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 59 32 0 data59x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 5 32 0 data5x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 60 32 0 data60x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 61 32 0 data61x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 62 32 0 data62x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 63 32 0 data63x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 6 32 0 data6x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 7 32 0 data7x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 8 32 0 data8x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 9 32 0 data9x 0 0 32 0
-- Retrieval info: CONNECT: @sel 0 0 6 0 sel 0 0 6 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL Chowdhury_LPM_32Bit64x1Mux_Dec7.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Chowdhury_LPM_32Bit64x1Mux_Dec7.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Chowdhury_LPM_32Bit64x1Mux_Dec7.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Chowdhury_LPM_32Bit64x1Mux_Dec7.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Chowdhury_LPM_32Bit64x1Mux_Dec7_inst.vhd FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Chowdhury_LPM_32Bit64x1Mux_Dec7_syn.v TRUE
-- Retrieval info: LIB_FILE: lpm
